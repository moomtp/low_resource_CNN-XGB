

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.types.all;

entity image_test is
    generic(TREE_RAM_BITS: positive := 14;
            NUM_CLASSES:   positive := 7;
            NUM_FEATURES:  positive := 35);
end image_test;

architecture behavior of image_test is
    
    component image
        generic(TREE_RAM_BITS: positive;
                NUM_CLASSES:   positive;
                NUM_FEATURES:  positive);
        port(-- Control signals
             Clk:   in std_logic;
             Reset: in std_logic;
             
             -- Inputs for the nodes reception (trees)
             Load_trees: in std_logic;
             Valid_node: in std_logic;
             Addr:       in std_logic_vector(TREE_RAM_BITS - 1  downto 0);
             Trees_din:  in std_logic_vector(31 downto 0);
             
             -- Inputs for the features reception (pixels)
             Load_features: in std_logic;
             Valid_feature: in std_logic;
             Features_din:  in std_logic_vector(15 downto 0);
             Last_feature:  in std_logic;
             
             -- Output signals
             --     Finish:     finish (also 'ready') signal
             --     Dout:       the selected class
             --     Greater:    the value of the selected class prediction
             --     Curr_state: the current state
             Finish:     out std_logic;
             Dout:       out std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);
             greater:    out std_logic_vector(31 downto 0);
             curr_state: out std_logic_vector(2 downto 0));
    end component;
    
    component counter is
        generic(BITS: natural);
        port(Clk:   in  std_logic;
             Reset: in  std_logic;
             Count: in  std_logic;
             Dout:  out std_logic_vector (BITS - 1 downto 0));
    end component;
    
    -- Inputs
    signal Clk:           std_logic := '0';
    signal Reset:         std_logic := '0';
    signal Load_trees:    std_logic := '0';
    signal Valid_node:    std_logic := '0';
    signal Addr:          std_logic_vector(TREE_RAM_BITS - 1 downto
                                           0) := (others => '0');
    signal Trees_din:     std_logic_vector(31 downto 0) := (others => '0');
    signal Load_features: std_logic := '0';
    signal Valid_feature: std_logic := '0';
    signal Features_din:  std_logic_vector(15 downto 0) := (others => '0');
    signal last_feature:  std_logic := '0';
    
    -- Outputs
    signal Finish:     std_logic;
    signal Dout:       std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);
    signal greater:    std_logic_vector(31 downto 0);
    signal curr_state: std_logic_vector(2 downto 0);
    
    -- Clock period definition
    constant Clk_period : time := 10 ns;
    
    -- Counter signals
    signal pc_count, hc_count: std_logic := '0';
    signal pixels, hits: std_logic_vector(15 downto 0) := (others => '0');
    
    -- Label signal
    signal class_label: std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);

begin
    
    -- Instantiate the Unit Under Test (UUT)
    uut: image
        generic map(TREE_RAM_BITS => TREE_RAM_BITS,
                    NUM_CLASSES   => NUM_CLASSES,
                    NUM_FEATURES  => NUM_FEATURES)
        port map(Clk           => Clk,
                 Reset         => Reset,
                 Load_trees    => Load_trees,
                 Valid_node    => Valid_node,
                 Addr          => Addr,
                 Trees_din     => Trees_din,
                 Load_features => Load_features,
                 Valid_feature => Valid_feature,
                 Features_din  => Features_din,
                 Last_feature  => Last_feature,
                 Finish        => Finish,
                 Dout          => Dout,
                 greater       => greater,
                 curr_state    => curr_state);
    
    -- To count the pixels
    pixel_counter: counter
        generic map(BITS => 16)
        port map(Clk   => Clk, 
                 Reset => Reset,
                 Count => pc_count,
                 Dout  => pixels);
    
    -- To count the hits
    hit_counter: counter
        generic map(BITS => 16)
        port map(Clk   => Clk, 
                 Reset => Reset,
                 Count => hc_count,
                 Dout  => hits);
    
    -- Clock process definition
    Clk_process: process
    begin
        Clk <= '0';
        wait for Clk_period/2;
        Clk <= '1';
        wait for Clk_period/2;
    end process;
    
    -- Stimulus process
    stim_proc: process
    begin
        
        Reset <= '1';
        
        -- hold reset state for 100 ns.
        wait for 100 ns;
        
        Reset <= '0';
        
        wait for Clk_period*10;
        


        
        -- LOAD TREES
        -----------------------------------------------------------------------
        
        -- Load and valid trees flags
        Load_trees <= '1';
        Valid_node <= '1';

        -- Class  0
        -----------
		Addr <=  "00000000000000";
		Trees_din <= x"010de978";
		wait for Clk_period;
		Addr <=  "00000000000001";
		Trees_din <= x"0108a438";
		wait for Clk_period;
		Addr <=  "00000000000010";
		Trees_din <= x"03fb9318";
		wait for Clk_period;
		Addr <=  "00000000000011";
		Trees_din <= x"0401a510";
		wait for Clk_period;
		Addr <=  "00000000000100";
		Trees_din <= x"1a013708";
		wait for Clk_period;
		Addr <=  "00000000000101";
		Trees_din <= x"0c000504";
		wait for Clk_period;
		Addr <=  "00000000000110";
		Trees_din <= x"ffab01ad";
		wait for Clk_period;
		Addr <=  "00000000000111";
		Trees_din <= x"ff5001ad";
		wait for Clk_period;
		Addr <=  "00000000001000";
		Trees_din <= x"0103d304";
		wait for Clk_period;
		Addr <=  "00000000001001";
		Trees_din <= x"ff8f01ad";
		wait for Clk_period;
		Addr <=  "00000000001010";
		Trees_din <= x"002701ad";
		wait for Clk_period;
		Addr <=  "00000000001011";
		Trees_din <= x"1c004104";
		wait for Clk_period;
		Addr <=  "00000000001100";
		Trees_din <= x"ff6601ad";
		wait for Clk_period;
		Addr <=  "00000000001101";
		Trees_din <= x"010b01ad";
		wait for Clk_period;
		Addr <=  "00000000001110";
		Trees_din <= x"0105bc10";
		wait for Clk_period;
		Addr <=  "00000000001111";
		Trees_din <= x"01017508";
		wait for Clk_period;
		Addr <=  "00000000010000";
		Trees_din <= x"1303b404";
		wait for Clk_period;
		Addr <=  "00000000010001";
		Trees_din <= x"ff5301ad";
		wait for Clk_period;
		Addr <=  "00000000010010";
		Trees_din <= x"000001ad";
		wait for Clk_period;
		Addr <=  "00000000010011";
		Trees_din <= x"1b002c04";
		wait for Clk_period;
		Addr <=  "00000000010100";
		Trees_din <= x"004101ad";
		wait for Clk_period;
		Addr <=  "00000000010101";
		Trees_din <= x"ff9301ad";
		wait for Clk_period;
		Addr <=  "00000000010110";
		Trees_din <= x"03000c08";
		wait for Clk_period;
		Addr <=  "00000000010111";
		Trees_din <= x"0afa1a04";
		wait for Clk_period;
		Addr <=  "00000000011000";
		Trees_din <= x"011f01ad";
		wait for Clk_period;
		Addr <=  "00000000011001";
		Trees_din <= x"ffd601ad";
		wait for Clk_period;
		Addr <=  "00000000011010";
		Trees_din <= x"1102eb04";
		wait for Clk_period;
		Addr <=  "00000000011011";
		Trees_din <= x"014801ad";
		wait for Clk_period;
		Addr <=  "00000000011100";
		Trees_din <= x"ff7001ad";
		wait for Clk_period;
		Addr <=  "00000000011101";
		Trees_din <= x"000f9e20";
		wait for Clk_period;
		Addr <=  "00000000011110";
		Trees_din <= x"02079810";
		wait for Clk_period;
		Addr <=  "00000000011111";
		Trees_din <= x"00090508";
		wait for Clk_period;
		Addr <=  "00000000100000";
		Trees_din <= x"040a4a04";
		wait for Clk_period;
		Addr <=  "00000000100001";
		Trees_din <= x"02b801ad";
		wait for Clk_period;
		Addr <=  "00000000100010";
		Trees_din <= x"005d01ad";
		wait for Clk_period;
		Addr <=  "00000000100011";
		Trees_din <= x"0400ad04";
		wait for Clk_period;
		Addr <=  "00000000100100";
		Trees_din <= x"01cd01ad";
		wait for Clk_period;
		Addr <=  "00000000100101";
		Trees_din <= x"ffb001ad";
		wait for Clk_period;
		Addr <=  "00000000100110";
		Trees_din <= x"18004d08";
		wait for Clk_period;
		Addr <=  "00000000100111";
		Trees_din <= x"0e02fe04";
		wait for Clk_period;
		Addr <=  "00000000101000";
		Trees_din <= x"ff9501ad";
		wait for Clk_period;
		Addr <=  "00000000101001";
		Trees_din <= x"00d401ad";
		wait for Clk_period;
		Addr <=  "00000000101010";
		Trees_din <= x"08006804";
		wait for Clk_period;
		Addr <=  "00000000101011";
		Trees_din <= x"ff9501ad";
		wait for Clk_period;
		Addr <=  "00000000101100";
		Trees_din <= x"025001ad";
		wait for Clk_period;
		Addr <=  "00000000101101";
		Trees_din <= x"0012ed10";
		wait for Clk_period;
		Addr <=  "00000000101110";
		Trees_din <= x"010c8d08";
		wait for Clk_period;
		Addr <=  "00000000101111";
		Trees_din <= x"05fbaf04";
		wait for Clk_period;
		Addr <=  "00000000110000";
		Trees_din <= x"ff8a01ad";
		wait for Clk_period;
		Addr <=  "00000000110001";
		Trees_din <= x"008a01ad";
		wait for Clk_period;
		Addr <=  "00000000110010";
		Trees_din <= x"04fb1404";
		wait for Clk_period;
		Addr <=  "00000000110011";
		Trees_din <= x"017101ad";
		wait for Clk_period;
		Addr <=  "00000000110100";
		Trees_din <= x"ffd001ad";
		wait for Clk_period;
		Addr <=  "00000000110101";
		Trees_din <= x"00164b08";
		wait for Clk_period;
		Addr <=  "00000000110110";
		Trees_din <= x"09005b04";
		wait for Clk_period;
		Addr <=  "00000000110111";
		Trees_din <= x"ff7901ad";
		wait for Clk_period;
		Addr <=  "00000000111000";
		Trees_din <= x"009d01ad";
		wait for Clk_period;
		Addr <=  "00000000111001";
		Trees_din <= x"1f000c04";
		wait for Clk_period;
		Addr <=  "00000000111010";
		Trees_din <= x"ff5001ad";
		wait for Clk_period;
		Addr <=  "00000000111011";
		Trees_din <= x"ffd001ad";
		wait for Clk_period;
		Addr <=  "00000000111100";
		Trees_din <= x"00100424";
		wait for Clk_period;
		Addr <=  "00000000111101";
		Trees_din <= x"020a7314";
		wait for Clk_period;
		Addr <=  "00000000111110";
		Trees_din <= x"01117e10";
		wait for Clk_period;
		Addr <=  "00000000111111";
		Trees_din <= x"03f97308";
		wait for Clk_period;
		Addr <=  "00000001000000";
		Trees_din <= x"17036004";
		wait for Clk_period;
		Addr <=  "00000001000001";
		Trees_din <= x"026001ad";
		wait for Clk_period;
		Addr <=  "00000001000010";
		Trees_din <= x"fff101ad";
		wait for Clk_period;
		Addr <=  "00000001000011";
		Trees_din <= x"11046104";
		wait for Clk_period;
		Addr <=  "00000001000100";
		Trees_din <= x"039801ad";
		wait for Clk_period;
		Addr <=  "00000001000101";
		Trees_din <= x"00b201ad";
		wait for Clk_period;
		Addr <=  "00000001000110";
		Trees_din <= x"03f701ad";
		wait for Clk_period;
		Addr <=  "00000001000111";
		Trees_din <= x"010fff08";
		wait for Clk_period;
		Addr <=  "00000001001000";
		Trees_din <= x"0008bf04";
		wait for Clk_period;
		Addr <=  "00000001001001";
		Trees_din <= x"00b201ad";
		wait for Clk_period;
		Addr <=  "00000001001010";
		Trees_din <= x"ff7301ad";
		wait for Clk_period;
		Addr <=  "00000001001011";
		Trees_din <= x"10028704";
		wait for Clk_period;
		Addr <=  "00000001001100";
		Trees_din <= x"024901ad";
		wait for Clk_period;
		Addr <=  "00000001001101";
		Trees_din <= x"ff9501ad";
		wait for Clk_period;
		Addr <=  "00000001001110";
		Trees_din <= x"0113e920";
		wait for Clk_period;
		Addr <=  "00000001001111";
		Trees_din <= x"00173a10";
		wait for Clk_period;
		Addr <=  "00000001010000";
		Trees_din <= x"0c02cf08";
		wait for Clk_period;
		Addr <=  "00000001010001";
		Trees_din <= x"0c001f04";
		wait for Clk_period;
		Addr <=  "00000001010010";
		Trees_din <= x"01c601ad";
		wait for Clk_period;
		Addr <=  "00000001010011";
		Trees_din <= x"ffff01ad";
		wait for Clk_period;
		Addr <=  "00000001010100";
		Trees_din <= x"18003c04";
		wait for Clk_period;
		Addr <=  "00000001010101";
		Trees_din <= x"fff701ad";
		wait for Clk_period;
		Addr <=  "00000001010110";
		Trees_din <= x"018701ad";
		wait for Clk_period;
		Addr <=  "00000001010111";
		Trees_din <= x"0112d608";
		wait for Clk_period;
		Addr <=  "00000001011000";
		Trees_din <= x"07004804";
		wait for Clk_period;
		Addr <=  "00000001011001";
		Trees_din <= x"003301ad";
		wait for Clk_period;
		Addr <=  "00000001011010";
		Trees_din <= x"ff5801ad";
		wait for Clk_period;
		Addr <=  "00000001011011";
		Trees_din <= x"01132a04";
		wait for Clk_period;
		Addr <=  "00000001011100";
		Trees_din <= x"00e201ad";
		wait for Clk_period;
		Addr <=  "00000001011101";
		Trees_din <= x"ff7501ad";
		wait for Clk_period;
		Addr <=  "00000001011110";
		Trees_din <= x"00161e0c";
		wait for Clk_period;
		Addr <=  "00000001011111";
		Trees_din <= x"1d005108";
		wait for Clk_period;
		Addr <=  "00000001100000";
		Trees_din <= x"11045104";
		wait for Clk_period;
		Addr <=  "00000001100001";
		Trees_din <= x"035e01ad";
		wait for Clk_period;
		Addr <=  "00000001100010";
		Trees_din <= x"00e201ad";
		wait for Clk_period;
		Addr <=  "00000001100011";
		Trees_din <= x"008e01ad";
		wait for Clk_period;
		Addr <=  "00000001100100";
		Trees_din <= x"01164208";
		wait for Clk_period;
		Addr <=  "00000001100101";
		Trees_din <= x"07005504";
		wait for Clk_period;
		Addr <=  "00000001100110";
		Trees_din <= x"002701ad";
		wait for Clk_period;
		Addr <=  "00000001100111";
		Trees_din <= x"ff6e01ad";
		wait for Clk_period;
		Addr <=  "00000001101000";
		Trees_din <= x"0801ca04";
		wait for Clk_period;
		Addr <=  "00000001101001";
		Trees_din <= x"002701ad";
		wait for Clk_period;
		Addr <=  "00000001101010";
		Trees_din <= x"01c601ad";
		wait for Clk_period;
		Addr <=  "00000001101011";
		Trees_din <= x"010cb458";
		wait for Clk_period;
		Addr <=  "00000001101100";
		Trees_din <= x"01084120";
		wait for Clk_period;
		Addr <=  "00000001101101";
		Trees_din <= x"000e0e1c";
		wait for Clk_period;
		Addr <=  "00000001101110";
		Trees_din <= x"0105bc10";
		wait for Clk_period;
		Addr <=  "00000001101111";
		Trees_din <= x"01017508";
		wait for Clk_period;
		Addr <=  "00000001110000";
		Trees_din <= x"1303b404";
		wait for Clk_period;
		Addr <=  "00000001110001";
		Trees_din <= x"ff5a0331";
		wait for Clk_period;
		Addr <=  "00000001110010";
		Trees_din <= x"000b0331";
		wait for Clk_period;
		Addr <=  "00000001110011";
		Trees_din <= x"1b002a04";
		wait for Clk_period;
		Addr <=  "00000001110100";
		Trees_din <= x"00510331";
		wait for Clk_period;
		Addr <=  "00000001110101";
		Trees_din <= x"ff9d0331";
		wait for Clk_period;
		Addr <=  "00000001110110";
		Trees_din <= x"020c6008";
		wait for Clk_period;
		Addr <=  "00000001110111";
		Trees_din <= x"07005c04";
		wait for Clk_period;
		Addr <=  "00000001111000";
		Trees_din <= x"00480331";
		wait for Clk_period;
		Addr <=  "00000001111001";
		Trees_din <= x"018e0331";
		wait for Clk_period;
		Addr <=  "00000001111010";
		Trees_din <= x"ff600331";
		wait for Clk_period;
		Addr <=  "00000001111011";
		Trees_din <= x"ff570331";
		wait for Clk_period;
		Addr <=  "00000001111100";
		Trees_din <= x"00100418";
		wait for Clk_period;
		Addr <=  "00000001111101";
		Trees_din <= x"0209130c";
		wait for Clk_period;
		Addr <=  "00000001111110";
		Trees_din <= x"1a008d04";
		wait for Clk_period;
		Addr <=  "00000001111111";
		Trees_din <= x"ff7a0331";
		wait for Clk_period;
		Addr <=  "00000010000000";
		Trees_din <= x"02022404";
		wait for Clk_period;
		Addr <=  "00000010000001";
		Trees_din <= x"01660331";
		wait for Clk_period;
		Addr <=  "00000010000010";
		Trees_din <= x"00c70331";
		wait for Clk_period;
		Addr <=  "00000010000011";
		Trees_din <= x"000e0e08";
		wait for Clk_period;
		Addr <=  "00000010000100";
		Trees_din <= x"09004c04";
		wait for Clk_period;
		Addr <=  "00000010000101";
		Trees_din <= x"00730331";
		wait for Clk_period;
		Addr <=  "00000010000110";
		Trees_din <= x"ff680331";
		wait for Clk_period;
		Addr <=  "00000010000111";
		Trees_din <= x"015e0331";
		wait for Clk_period;
		Addr <=  "00000010001000";
		Trees_din <= x"00153210";
		wait for Clk_period;
		Addr <=  "00000010001001";
		Trees_din <= x"0c028608";
		wait for Clk_period;
		Addr <=  "00000010001010";
		Trees_din <= x"1603fe04";
		wait for Clk_period;
		Addr <=  "00000010001011";
		Trees_din <= x"ff660331";
		wait for Clk_period;
		Addr <=  "00000010001100";
		Trees_din <= x"00860331";
		wait for Clk_period;
		Addr <=  "00000010001101";
		Trees_din <= x"0bfa1604";
		wait for Clk_period;
		Addr <=  "00000010001110";
		Trees_din <= x"01020331";
		wait for Clk_period;
		Addr <=  "00000010001111";
		Trees_din <= x"ffbc0331";
		wait for Clk_period;
		Addr <=  "00000010010000";
		Trees_din <= x"1f000c08";
		wait for Clk_period;
		Addr <=  "00000010010001";
		Trees_din <= x"03f88c04";
		wait for Clk_period;
		Addr <=  "00000010010010";
		Trees_din <= x"ff560331";
		wait for Clk_period;
		Addr <=  "00000010010011";
		Trees_din <= x"ffc40331";
		wait for Clk_period;
		Addr <=  "00000010010100";
		Trees_din <= x"0b03cc04";
		wait for Clk_period;
		Addr <=  "00000010010101";
		Trees_din <= x"ffa00331";
		wait for Clk_period;
		Addr <=  "00000010010110";
		Trees_din <= x"00420331";
		wait for Clk_period;
		Addr <=  "00000010010111";
		Trees_din <= x"00138a30";
		wait for Clk_period;
		Addr <=  "00000010011000";
		Trees_din <= x"020baf20";
		wait for Clk_period;
		Addr <=  "00000010011001";
		Trees_din <= x"010f7410";
		wait for Clk_period;
		Addr <=  "00000010011010";
		Trees_din <= x"000f3608";
		wait for Clk_period;
		Addr <=  "00000010011011";
		Trees_din <= x"14001804";
		wait for Clk_period;
		Addr <=  "00000010011100";
		Trees_din <= x"ffc50331";
		wait for Clk_period;
		Addr <=  "00000010011101";
		Trees_din <= x"01620331";
		wait for Clk_period;
		Addr <=  "00000010011110";
		Trees_din <= x"0bfa2304";
		wait for Clk_period;
		Addr <=  "00000010011111";
		Trees_din <= x"ff9a0331";
		wait for Clk_period;
		Addr <=  "00000010100000";
		Trees_din <= x"00a00331";
		wait for Clk_period;
		Addr <=  "00000010100001";
		Trees_din <= x"22000008";
		wait for Clk_period;
		Addr <=  "00000010100010";
		Trees_din <= x"0113e904";
		wait for Clk_period;
		Addr <=  "00000010100011";
		Trees_din <= x"01790331";
		wait for Clk_period;
		Addr <=  "00000010100100";
		Trees_din <= x"01ba0331";
		wait for Clk_period;
		Addr <=  "00000010100101";
		Trees_din <= x"17002104";
		wait for Clk_period;
		Addr <=  "00000010100110";
		Trees_din <= x"ff8f0331";
		wait for Clk_period;
		Addr <=  "00000010100111";
		Trees_din <= x"012b0331";
		wait for Clk_period;
		Addr <=  "00000010101000";
		Trees_din <= x"17000908";
		wait for Clk_period;
		Addr <=  "00000010101001";
		Trees_din <= x"0c01bf04";
		wait for Clk_period;
		Addr <=  "00000010101010";
		Trees_din <= x"00260331";
		wait for Clk_period;
		Addr <=  "00000010101011";
		Trees_din <= x"01520331";
		wait for Clk_period;
		Addr <=  "00000010101100";
		Trees_din <= x"10fad204";
		wait for Clk_period;
		Addr <=  "00000010101101";
		Trees_din <= x"00b20331";
		wait for Clk_period;
		Addr <=  "00000010101110";
		Trees_din <= x"ff660331";
		wait for Clk_period;
		Addr <=  "00000010101111";
		Trees_din <= x"01128f20";
		wait for Clk_period;
		Addr <=  "00000010110000";
		Trees_din <= x"0017f910";
		wait for Clk_period;
		Addr <=  "00000010110001";
		Trees_din <= x"1402ad08";
		wait for Clk_period;
		Addr <=  "00000010110010";
		Trees_din <= x"0f000004";
		wait for Clk_period;
		Addr <=  "00000010110011";
		Trees_din <= x"00be0331";
		wait for Clk_period;
		Addr <=  "00000010110100";
		Trees_din <= x"ff880331";
		wait for Clk_period;
		Addr <=  "00000010110101";
		Trees_din <= x"010ea204";
		wait for Clk_period;
		Addr <=  "00000010110110";
		Trees_din <= x"ffde0331";
		wait for Clk_period;
		Addr <=  "00000010110111";
		Trees_din <= x"01050331";
		wait for Clk_period;
		Addr <=  "00000010111000";
		Trees_din <= x"18004f08";
		wait for Clk_period;
		Addr <=  "00000010111001";
		Trees_din <= x"03f53b04";
		wait for Clk_period;
		Addr <=  "00000010111010";
		Trees_din <= x"ff580331";
		wait for Clk_period;
		Addr <=  "00000010111011";
		Trees_din <= x"ffc40331";
		wait for Clk_period;
		Addr <=  "00000010111100";
		Trees_din <= x"07005604";
		wait for Clk_period;
		Addr <=  "00000010111101";
		Trees_din <= x"00bc0331";
		wait for Clk_period;
		Addr <=  "00000010111110";
		Trees_din <= x"ff8b0331";
		wait for Clk_period;
		Addr <=  "00000010111111";
		Trees_din <= x"0018d010";
		wait for Clk_period;
		Addr <=  "00000011000000";
		Trees_din <= x"13012a08";
		wait for Clk_period;
		Addr <=  "00000011000001";
		Trees_din <= x"0d023e04";
		wait for Clk_period;
		Addr <=  "00000011000010";
		Trees_din <= x"019b0331";
		wait for Clk_period;
		Addr <=  "00000011000011";
		Trees_din <= x"00650331";
		wait for Clk_period;
		Addr <=  "00000011000100";
		Trees_din <= x"17000004";
		wait for Clk_period;
		Addr <=  "00000011000101";
		Trees_din <= x"00360331";
		wait for Clk_period;
		Addr <=  "00000011000110";
		Trees_din <= x"ff860331";
		wait for Clk_period;
		Addr <=  "00000011000111";
		Trees_din <= x"0c02cf04";
		wait for Clk_period;
		Addr <=  "00000011001000";
		Trees_din <= x"ff660331";
		wait for Clk_period;
		Addr <=  "00000011001001";
		Trees_din <= x"0c036404";
		wait for Clk_period;
		Addr <=  "00000011001010";
		Trees_din <= x"016e0331";
		wait for Clk_period;
		Addr <=  "00000011001011";
		Trees_din <= x"ffa50331";
		wait for Clk_period;
		Addr <=  "00000011001100";
		Trees_din <= x"010b116c";
		wait for Clk_period;
		Addr <=  "00000011001101";
		Trees_din <= x"0105bc34";
		wait for Clk_period;
		Addr <=  "00000011001110";
		Trees_din <= x"03fc9714";
		wait for Clk_period;
		Addr <=  "00000011001111";
		Trees_din <= x"0af74908";
		wait for Clk_period;
		Addr <=  "00000011010000";
		Trees_din <= x"09005504";
		wait for Clk_period;
		Addr <=  "00000011010001";
		Trees_din <= x"003704d5";
		wait for Clk_period;
		Addr <=  "00000011010010";
		Trees_din <= x"ffa304d5";
		wait for Clk_period;
		Addr <=  "00000011010011";
		Trees_din <= x"0105aa04";
		wait for Clk_period;
		Addr <=  "00000011010100";
		Trees_din <= x"ff5904d5";
		wait for Clk_period;
		Addr <=  "00000011010101";
		Trees_din <= x"1a00ce04";
		wait for Clk_period;
		Addr <=  "00000011010110";
		Trees_din <= x"003d04d5";
		wait for Clk_period;
		Addr <=  "00000011010111";
		Trees_din <= x"ff9404d5";
		wait for Clk_period;
		Addr <=  "00000011011000";
		Trees_din <= x"01017510";
		wait for Clk_period;
		Addr <=  "00000011011001";
		Trees_din <= x"0f03e608";
		wait for Clk_period;
		Addr <=  "00000011011010";
		Trees_din <= x"03fce704";
		wait for Clk_period;
		Addr <=  "00000011011011";
		Trees_din <= x"ffdf04d5";
		wait for Clk_period;
		Addr <=  "00000011011100";
		Trees_din <= x"ff5a04d5";
		wait for Clk_period;
		Addr <=  "00000011011101";
		Trees_din <= x"16005204";
		wait for Clk_period;
		Addr <=  "00000011011110";
		Trees_din <= x"ff8904d5";
		wait for Clk_period;
		Addr <=  "00000011011111";
		Trees_din <= x"00e004d5";
		wait for Clk_period;
		Addr <=  "00000011100000";
		Trees_din <= x"0d019308";
		wait for Clk_period;
		Addr <=  "00000011100001";
		Trees_din <= x"06fcc204";
		wait for Clk_period;
		Addr <=  "00000011100010";
		Trees_din <= x"ff7a04d5";
		wait for Clk_period;
		Addr <=  "00000011100011";
		Trees_din <= x"003904d5";
		wait for Clk_period;
		Addr <=  "00000011100100";
		Trees_din <= x"13ffd004";
		wait for Clk_period;
		Addr <=  "00000011100101";
		Trees_din <= x"ffd204d5";
		wait for Clk_period;
		Addr <=  "00000011100110";
		Trees_din <= x"007b04d5";
		wait for Clk_period;
		Addr <=  "00000011100111";
		Trees_din <= x"0010b120";
		wait for Clk_period;
		Addr <=  "00000011101000";
		Trees_din <= x"020baf10";
		wait for Clk_period;
		Addr <=  "00000011101001";
		Trees_din <= x"0ef9de08";
		wait for Clk_period;
		Addr <=  "00000011101010";
		Trees_din <= x"00060104";
		wait for Clk_period;
		Addr <=  "00000011101011";
		Trees_din <= x"01b804d5";
		wait for Clk_period;
		Addr <=  "00000011101100";
		Trees_din <= x"004504d5";
		wait for Clk_period;
		Addr <=  "00000011101101";
		Trees_din <= x"0202f304";
		wait for Clk_period;
		Addr <=  "00000011101110";
		Trees_din <= x"008d04d5";
		wait for Clk_period;
		Addr <=  "00000011101111";
		Trees_din <= x"000d04d5";
		wait for Clk_period;
		Addr <=  "00000011110000";
		Trees_din <= x"09004f08";
		wait for Clk_period;
		Addr <=  "00000011110001";
		Trees_din <= x"10020304";
		wait for Clk_period;
		Addr <=  "00000011110010";
		Trees_din <= x"00c804d5";
		wait for Clk_period;
		Addr <=  "00000011110011";
		Trees_din <= x"ff7b04d5";
		wait for Clk_period;
		Addr <=  "00000011110100";
		Trees_din <= x"0009b104";
		wait for Clk_period;
		Addr <=  "00000011110101";
		Trees_din <= x"ff6204d5";
		wait for Clk_period;
		Addr <=  "00000011110110";
		Trees_din <= x"ffed04d5";
		wait for Clk_period;
		Addr <=  "00000011110111";
		Trees_din <= x"0014d00c";
		wait for Clk_period;
		Addr <=  "00000011111000";
		Trees_din <= x"0a044c08";
		wait for Clk_period;
		Addr <=  "00000011111001";
		Trees_din <= x"0af89204";
		wait for Clk_period;
		Addr <=  "00000011111010";
		Trees_din <= x"004004d5";
		wait for Clk_period;
		Addr <=  "00000011111011";
		Trees_din <= x"ff7e04d5";
		wait for Clk_period;
		Addr <=  "00000011111100";
		Trees_din <= x"009704d5";
		wait for Clk_period;
		Addr <=  "00000011111101";
		Trees_din <= x"03fa9f08";
		wait for Clk_period;
		Addr <=  "00000011111110";
		Trees_din <= x"21000004";
		wait for Clk_period;
		Addr <=  "00000011111111";
		Trees_din <= x"ff5a04d5";
		wait for Clk_period;
		Addr <=  "00000100000000";
		Trees_din <= x"ffa004d5";
		wait for Clk_period;
		Addr <=  "00000100000001";
		Trees_din <= x"001e04d5";
		wait for Clk_period;
		Addr <=  "00000100000010";
		Trees_din <= x"00138a38";
		wait for Clk_period;
		Addr <=  "00000100000011";
		Trees_din <= x"010f7420";
		wait for Clk_period;
		Addr <=  "00000100000100";
		Trees_din <= x"020b0110";
		wait for Clk_period;
		Addr <=  "00000100000101";
		Trees_din <= x"000f6f08";
		wait for Clk_period;
		Addr <=  "00000100000110";
		Trees_din <= x"02011804";
		wait for Clk_period;
		Addr <=  "00000100000111";
		Trees_din <= x"013e04d5";
		wait for Clk_period;
		Addr <=  "00000100001000";
		Trees_din <= x"00b404d5";
		wait for Clk_period;
		Addr <=  "00000100001001";
		Trees_din <= x"05fbaf04";
		wait for Clk_period;
		Addr <=  "00000100001010";
		Trees_din <= x"001e04d5";
		wait for Clk_period;
		Addr <=  "00000100001011";
		Trees_din <= x"015f04d5";
		wait for Clk_period;
		Addr <=  "00000100001100";
		Trees_din <= x"0c02ae08";
		wait for Clk_period;
		Addr <=  "00000100001101";
		Trees_din <= x"05fb4104";
		wait for Clk_period;
		Addr <=  "00000100001110";
		Trees_din <= x"ff6604d5";
		wait for Clk_period;
		Addr <=  "00000100001111";
		Trees_din <= x"003a04d5";
		wait for Clk_period;
		Addr <=  "00000100010000";
		Trees_din <= x"00079004";
		wait for Clk_period;
		Addr <=  "00000100010001";
		Trees_din <= x"013404d5";
		wait for Clk_period;
		Addr <=  "00000100010010";
		Trees_din <= x"ffa004d5";
		wait for Clk_period;
		Addr <=  "00000100010011";
		Trees_din <= x"000fd30c";
		wait for Clk_period;
		Addr <=  "00000100010100";
		Trees_din <= x"15007104";
		wait for Clk_period;
		Addr <=  "00000100010101";
		Trees_din <= x"002504d5";
		wait for Clk_period;
		Addr <=  "00000100010110";
		Trees_din <= x"020a7304";
		wait for Clk_period;
		Addr <=  "00000100010111";
		Trees_din <= x"012a04d5";
		wait for Clk_period;
		Addr <=  "00000100011000";
		Trees_din <= x"008c04d5";
		wait for Clk_period;
		Addr <=  "00000100011001";
		Trees_din <= x"0efb2404";
		wait for Clk_period;
		Addr <=  "00000100011010";
		Trees_din <= x"ff7104d5";
		wait for Clk_period;
		Addr <=  "00000100011011";
		Trees_din <= x"1c004304";
		wait for Clk_period;
		Addr <=  "00000100011100";
		Trees_din <= x"010a04d5";
		wait for Clk_period;
		Addr <=  "00000100011101";
		Trees_din <= x"002904d5";
		wait for Clk_period;
		Addr <=  "00000100011110";
		Trees_din <= x"01128f18";
		wait for Clk_period;
		Addr <=  "00000100011111";
		Trees_din <= x"0015320c";
		wait for Clk_period;
		Addr <=  "00000100100000";
		Trees_din <= x"0d029108";
		wait for Clk_period;
		Addr <=  "00000100100001";
		Trees_din <= x"00146004";
		wait for Clk_period;
		Addr <=  "00000100100010";
		Trees_din <= x"ff7504d5";
		wait for Clk_period;
		Addr <=  "00000100100011";
		Trees_din <= x"010b04d5";
		wait for Clk_period;
		Addr <=  "00000100100100";
		Trees_din <= x"ff6c04d5";
		wait for Clk_period;
		Addr <=  "00000100100101";
		Trees_din <= x"21000308";
		wait for Clk_period;
		Addr <=  "00000100100110";
		Trees_din <= x"03f7f004";
		wait for Clk_period;
		Addr <=  "00000100100111";
		Trees_din <= x"ff6d04d5";
		wait for Clk_period;
		Addr <=  "00000100101000";
		Trees_din <= x"002f04d5";
		wait for Clk_period;
		Addr <=  "00000100101001";
		Trees_din <= x"007804d5";
		wait for Clk_period;
		Addr <=  "00000100101010";
		Trees_din <= x"001ac110";
		wait for Clk_period;
		Addr <=  "00000100101011";
		Trees_din <= x"13012a08";
		wait for Clk_period;
		Addr <=  "00000100101100";
		Trees_din <= x"1d004f04";
		wait for Clk_period;
		Addr <=  "00000100101101";
		Trees_din <= x"010004d5";
		wait for Clk_period;
		Addr <=  "00000100101110";
		Trees_din <= x"ffd404d5";
		wait for Clk_period;
		Addr <=  "00000100101111";
		Trees_din <= x"0bfae904";
		wait for Clk_period;
		Addr <=  "00000100110000";
		Trees_din <= x"003a04d5";
		wait for Clk_period;
		Addr <=  "00000100110001";
		Trees_din <= x"ff8504d5";
		wait for Clk_period;
		Addr <=  "00000100110010";
		Trees_din <= x"10fb4004";
		wait for Clk_period;
		Addr <=  "00000100110011";
		Trees_din <= x"007f04d5";
		wait for Clk_period;
		Addr <=  "00000100110100";
		Trees_din <= x"ff7004d5";
		wait for Clk_period;
		Addr <=  "00000100110101";
		Trees_din <= x"010b1164";
		wait for Clk_period;
		Addr <=  "00000100110110";
		Trees_din <= x"0010b13c";
		wait for Clk_period;
		Addr <=  "00000100110111";
		Trees_din <= x"0105bc20";
		wait for Clk_period;
		Addr <=  "00000100111000";
		Trees_din <= x"01017510";
		wait for Clk_period;
		Addr <=  "00000100111001";
		Trees_din <= x"1303b408";
		wait for Clk_period;
		Addr <=  "00000100111010";
		Trees_din <= x"09005e04";
		wait for Clk_period;
		Addr <=  "00000100111011";
		Trees_din <= x"ff610669";
		wait for Clk_period;
		Addr <=  "00000100111100";
		Trees_din <= x"fff30669";
		wait for Clk_period;
		Addr <=  "00000100111101";
		Trees_din <= x"19008904";
		wait for Clk_period;
		Addr <=  "00000100111110";
		Trees_din <= x"00d40669";
		wait for Clk_period;
		Addr <=  "00000100111111";
		Trees_din <= x"ff920669";
		wait for Clk_period;
		Addr <=  "00000101000000";
		Trees_din <= x"03fc9708";
		wait for Clk_period;
		Addr <=  "00000101000001";
		Trees_din <= x"18005304";
		wait for Clk_period;
		Addr <=  "00000101000010";
		Trees_din <= x"ff5f0669";
		wait for Clk_period;
		Addr <=  "00000101000011";
		Trees_din <= x"00330669";
		wait for Clk_period;
		Addr <=  "00000101000100";
		Trees_din <= x"0d019304";
		wait for Clk_period;
		Addr <=  "00000101000101";
		Trees_din <= x"ff9c0669";
		wait for Clk_period;
		Addr <=  "00000101000110";
		Trees_din <= x"001d0669";
		wait for Clk_period;
		Addr <=  "00000101000111";
		Trees_din <= x"020d0610";
		wait for Clk_period;
		Addr <=  "00000101001000";
		Trees_din <= x"13014108";
		wait for Clk_period;
		Addr <=  "00000101001001";
		Trees_din <= x"06f61f04";
		wait for Clk_period;
		Addr <=  "00000101001010";
		Trees_din <= x"003c0669";
		wait for Clk_period;
		Addr <=  "00000101001011";
		Trees_din <= x"00a30669";
		wait for Clk_period;
		Addr <=  "00000101001100";
		Trees_din <= x"11fcaf04";
		wait for Clk_period;
		Addr <=  "00000101001101";
		Trees_din <= x"00dc0669";
		wait for Clk_period;
		Addr <=  "00000101001110";
		Trees_din <= x"ffab0669";
		wait for Clk_period;
		Addr <=  "00000101001111";
		Trees_din <= x"0e03b208";
		wait for Clk_period;
		Addr <=  "00000101010000";
		Trees_din <= x"18004b04";
		wait for Clk_period;
		Addr <=  "00000101010001";
		Trees_din <= x"ff660669";
		wait for Clk_period;
		Addr <=  "00000101010010";
		Trees_din <= x"00360669";
		wait for Clk_period;
		Addr <=  "00000101010011";
		Trees_din <= x"007f0669";
		wait for Clk_period;
		Addr <=  "00000101010100";
		Trees_din <= x"0014d014";
		wait for Clk_period;
		Addr <=  "00000101010101";
		Trees_din <= x"0105aa04";
		wait for Clk_period;
		Addr <=  "00000101010110";
		Trees_din <= x"ff600669";
		wait for Clk_period;
		Addr <=  "00000101010111";
		Trees_din <= x"0012ed08";
		wait for Clk_period;
		Addr <=  "00000101011000";
		Trees_din <= x"14001b04";
		wait for Clk_period;
		Addr <=  "00000101011001";
		Trees_din <= x"00300669";
		wait for Clk_period;
		Addr <=  "00000101011010";
		Trees_din <= x"ff640669";
		wait for Clk_period;
		Addr <=  "00000101011011";
		Trees_din <= x"06f5a604";
		wait for Clk_period;
		Addr <=  "00000101011100";
		Trees_din <= x"ff750669";
		wait for Clk_period;
		Addr <=  "00000101011101";
		Trees_din <= x"00760669";
		wait for Clk_period;
		Addr <=  "00000101011110";
		Trees_din <= x"03faba0c";
		wait for Clk_period;
		Addr <=  "00000101011111";
		Trees_din <= x"0d000008";
		wait for Clk_period;
		Addr <=  "00000101100000";
		Trees_din <= x"1a00dd04";
		wait for Clk_period;
		Addr <=  "00000101100001";
		Trees_din <= x"ff740669";
		wait for Clk_period;
		Addr <=  "00000101100010";
		Trees_din <= x"003e0669";
		wait for Clk_period;
		Addr <=  "00000101100011";
		Trees_din <= x"ff5d0669";
		wait for Clk_period;
		Addr <=  "00000101100100";
		Trees_din <= x"05f93f04";
		wait for Clk_period;
		Addr <=  "00000101100101";
		Trees_din <= x"00450669";
		wait for Clk_period;
		Addr <=  "00000101100110";
		Trees_din <= x"ff770669";
		wait for Clk_period;
		Addr <=  "00000101100111";
		Trees_din <= x"0015323c";
		wait for Clk_period;
		Addr <=  "00000101101000";
		Trees_din <= x"01114420";
		wait for Clk_period;
		Addr <=  "00000101101001";
		Trees_din <= x"00115710";
		wait for Clk_period;
		Addr <=  "00000101101010";
		Trees_din <= x"020b0108";
		wait for Clk_period;
		Addr <=  "00000101101011";
		Trees_din <= x"06f65504";
		wait for Clk_period;
		Addr <=  "00000101101100";
		Trees_din <= x"00980669";
		wait for Clk_period;
		Addr <=  "00000101101101";
		Trees_din <= x"00e90669";
		wait for Clk_period;
		Addr <=  "00000101101110";
		Trees_din <= x"1c003604";
		wait for Clk_period;
		Addr <=  "00000101101111";
		Trees_din <= x"ff8a0669";
		wait for Clk_period;
		Addr <=  "00000101110000";
		Trees_din <= x"007d0669";
		wait for Clk_period;
		Addr <=  "00000101110001";
		Trees_din <= x"05fbaf08";
		wait for Clk_period;
		Addr <=  "00000101110010";
		Trees_din <= x"010cb404";
		wait for Clk_period;
		Addr <=  "00000101110011";
		Trees_din <= x"ff690669";
		wait for Clk_period;
		Addr <=  "00000101110100";
		Trees_din <= x"00180669";
		wait for Clk_period;
		Addr <=  "00000101110101";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00000101110110";
		Trees_din <= x"ff9e0669";
		wait for Clk_period;
		Addr <=  "00000101110111";
		Trees_din <= x"01670669";
		wait for Clk_period;
		Addr <=  "00000101111000";
		Trees_din <= x"0113e910";
		wait for Clk_period;
		Addr <=  "00000101111001";
		Trees_din <= x"0afccc08";
		wait for Clk_period;
		Addr <=  "00000101111010";
		Trees_din <= x"08000004";
		wait for Clk_period;
		Addr <=  "00000101111011";
		Trees_din <= x"000b0669";
		wait for Clk_period;
		Addr <=  "00000101111100";
		Trees_din <= x"00fc0669";
		wait for Clk_period;
		Addr <=  "00000101111101";
		Trees_din <= x"0f000c04";
		wait for Clk_period;
		Addr <=  "00000101111110";
		Trees_din <= x"ff770669";
		wait for Clk_period;
		Addr <=  "00000101111111";
		Trees_din <= x"009b0669";
		wait for Clk_period;
		Addr <=  "00000110000000";
		Trees_din <= x"22000008";
		wait for Clk_period;
		Addr <=  "00000110000001";
		Trees_din <= x"07004904";
		wait for Clk_period;
		Addr <=  "00000110000010";
		Trees_din <= x"00500669";
		wait for Clk_period;
		Addr <=  "00000110000011";
		Trees_din <= x"01010669";
		wait for Clk_period;
		Addr <=  "00000110000100";
		Trees_din <= x"00080669";
		wait for Clk_period;
		Addr <=  "00000110000101";
		Trees_din <= x"01128f14";
		wait for Clk_period;
		Addr <=  "00000110000110";
		Trees_din <= x"21000310";
		wait for Clk_period;
		Addr <=  "00000110000111";
		Trees_din <= x"07004808";
		wait for Clk_period;
		Addr <=  "00000110001000";
		Trees_din <= x"0a02b704";
		wait for Clk_period;
		Addr <=  "00000110001001";
		Trees_din <= x"ffa40669";
		wait for Clk_period;
		Addr <=  "00000110001010";
		Trees_din <= x"00de0669";
		wait for Clk_period;
		Addr <=  "00000110001011";
		Trees_din <= x"0bf74e04";
		wait for Clk_period;
		Addr <=  "00000110001100";
		Trees_din <= x"003b0669";
		wait for Clk_period;
		Addr <=  "00000110001101";
		Trees_din <= x"ff710669";
		wait for Clk_period;
		Addr <=  "00000110001110";
		Trees_din <= x"00750669";
		wait for Clk_period;
		Addr <=  "00000110001111";
		Trees_din <= x"11ffce08";
		wait for Clk_period;
		Addr <=  "00000110010000";
		Trees_din <= x"01164204";
		wait for Clk_period;
		Addr <=  "00000110010001";
		Trees_din <= x"ff780669";
		wait for Clk_period;
		Addr <=  "00000110010010";
		Trees_din <= x"00290669";
		wait for Clk_period;
		Addr <=  "00000110010011";
		Trees_din <= x"0f02a808";
		wait for Clk_period;
		Addr <=  "00000110010100";
		Trees_din <= x"1c002904";
		wait for Clk_period;
		Addr <=  "00000110010101";
		Trees_din <= x"ff910669";
		wait for Clk_period;
		Addr <=  "00000110010110";
		Trees_din <= x"00e60669";
		wait for Clk_period;
		Addr <=  "00000110010111";
		Trees_din <= x"05f77304";
		wait for Clk_period;
		Addr <=  "00000110011000";
		Trees_din <= x"00300669";
		wait for Clk_period;
		Addr <=  "00000110011001";
		Trees_din <= x"ff7f0669";
		wait for Clk_period;
		Addr <=  "00000110011010";
		Trees_din <= x"0108a460";
		wait for Clk_period;
		Addr <=  "00000110011011";
		Trees_din <= x"03fa9f28";
		wait for Clk_period;
		Addr <=  "00000110011100";
		Trees_din <= x"03f87814";
		wait for Clk_period;
		Addr <=  "00000110011101";
		Trees_din <= x"04fe5b0c";
		wait for Clk_period;
		Addr <=  "00000110011110";
		Trees_din <= x"0d000008";
		wait for Clk_period;
		Addr <=  "00000110011111";
		Trees_din <= x"15009c04";
		wait for Clk_period;
		Addr <=  "00000110100000";
		Trees_din <= x"ff7d07fd";
		wait for Clk_period;
		Addr <=  "00000110100001";
		Trees_din <= x"003907fd";
		wait for Clk_period;
		Addr <=  "00000110100010";
		Trees_din <= x"ff6007fd";
		wait for Clk_period;
		Addr <=  "00000110100011";
		Trees_din <= x"14019f04";
		wait for Clk_period;
		Addr <=  "00000110100100";
		Trees_din <= x"004507fd";
		wait for Clk_period;
		Addr <=  "00000110100101";
		Trees_din <= x"ff9d07fd";
		wait for Clk_period;
		Addr <=  "00000110100110";
		Trees_din <= x"03f9110c";
		wait for Clk_period;
		Addr <=  "00000110100111";
		Trees_din <= x"0105aa04";
		wait for Clk_period;
		Addr <=  "00000110101000";
		Trees_din <= x"ff6b07fd";
		wait for Clk_period;
		Addr <=  "00000110101001";
		Trees_din <= x"0106e504";
		wait for Clk_period;
		Addr <=  "00000110101010";
		Trees_din <= x"016907fd";
		wait for Clk_period;
		Addr <=  "00000110101011";
		Trees_din <= x"ffd807fd";
		wait for Clk_period;
		Addr <=  "00000110101100";
		Trees_din <= x"07005e04";
		wait for Clk_period;
		Addr <=  "00000110101101";
		Trees_din <= x"ff6007fd";
		wait for Clk_period;
		Addr <=  "00000110101110";
		Trees_din <= x"002907fd";
		wait for Clk_period;
		Addr <=  "00000110101111";
		Trees_din <= x"01017518";
		wait for Clk_period;
		Addr <=  "00000110110000";
		Trees_din <= x"0f03e60c";
		wait for Clk_period;
		Addr <=  "00000110110001";
		Trees_din <= x"07005e04";
		wait for Clk_period;
		Addr <=  "00000110110010";
		Trees_din <= x"ff6007fd";
		wait for Clk_period;
		Addr <=  "00000110110011";
		Trees_din <= x"0f003004";
		wait for Clk_period;
		Addr <=  "00000110110100";
		Trees_din <= x"ffa507fd";
		wait for Clk_period;
		Addr <=  "00000110110101";
		Trees_din <= x"004707fd";
		wait for Clk_period;
		Addr <=  "00000110110110";
		Trees_din <= x"16005208";
		wait for Clk_period;
		Addr <=  "00000110110111";
		Trees_din <= x"12fe6204";
		wait for Clk_period;
		Addr <=  "00000110111000";
		Trees_din <= x"003507fd";
		wait for Clk_period;
		Addr <=  "00000110111001";
		Trees_din <= x"ff7407fd";
		wait for Clk_period;
		Addr <=  "00000110111010";
		Trees_din <= x"00b907fd";
		wait for Clk_period;
		Addr <=  "00000110111011";
		Trees_din <= x"0105bc10";
		wait for Clk_period;
		Addr <=  "00000110111100";
		Trees_din <= x"0d019308";
		wait for Clk_period;
		Addr <=  "00000110111101";
		Trees_din <= x"06fcc204";
		wait for Clk_period;
		Addr <=  "00000110111110";
		Trees_din <= x"ff8307fd";
		wait for Clk_period;
		Addr <=  "00000110111111";
		Trees_din <= x"003e07fd";
		wait for Clk_period;
		Addr <=  "00000111000000";
		Trees_din <= x"0d020204";
		wait for Clk_period;
		Addr <=  "00000111000001";
		Trees_din <= x"008c07fd";
		wait for Clk_period;
		Addr <=  "00000111000010";
		Trees_din <= x"ffda07fd";
		wait for Clk_period;
		Addr <=  "00000111000011";
		Trees_din <= x"15009908";
		wait for Clk_period;
		Addr <=  "00000111000100";
		Trees_din <= x"11032704";
		wait for Clk_period;
		Addr <=  "00000111000101";
		Trees_din <= x"009007fd";
		wait for Clk_period;
		Addr <=  "00000111000110";
		Trees_din <= x"ff7107fd";
		wait for Clk_period;
		Addr <=  "00000111000111";
		Trees_din <= x"18003c04";
		wait for Clk_period;
		Addr <=  "00000111001000";
		Trees_din <= x"002b07fd";
		wait for Clk_period;
		Addr <=  "00000111001001";
		Trees_din <= x"ff7707fd";
		wait for Clk_period;
		Addr <=  "00000111001010";
		Trees_din <= x"00167640";
		wait for Clk_period;
		Addr <=  "00000111001011";
		Trees_din <= x"010f7420";
		wait for Clk_period;
		Addr <=  "00000111001100";
		Trees_din <= x"0011cf10";
		wait for Clk_period;
		Addr <=  "00000111001101";
		Trees_din <= x"020b0108";
		wait for Clk_period;
		Addr <=  "00000111001110";
		Trees_din <= x"09005d04";
		wait for Clk_period;
		Addr <=  "00000111001111";
		Trees_din <= x"007d07fd";
		wait for Clk_period;
		Addr <=  "00000111010000";
		Trees_din <= x"ff7d07fd";
		wait for Clk_period;
		Addr <=  "00000111010001";
		Trees_din <= x"0e045004";
		wait for Clk_period;
		Addr <=  "00000111010010";
		Trees_din <= x"ffb407fd";
		wait for Clk_period;
		Addr <=  "00000111010011";
		Trees_din <= x"014d07fd";
		wait for Clk_period;
		Addr <=  "00000111010100";
		Trees_din <= x"08015b08";
		wait for Clk_period;
		Addr <=  "00000111010101";
		Trees_din <= x"0e03d004";
		wait for Clk_period;
		Addr <=  "00000111010110";
		Trees_din <= x"ff8407fd";
		wait for Clk_period;
		Addr <=  "00000111010111";
		Trees_din <= x"00ab07fd";
		wait for Clk_period;
		Addr <=  "00000111011000";
		Trees_din <= x"15009804";
		wait for Clk_period;
		Addr <=  "00000111011001";
		Trees_din <= x"ffbc07fd";
		wait for Clk_period;
		Addr <=  "00000111011010";
		Trees_din <= x"00cc07fd";
		wait for Clk_period;
		Addr <=  "00000111011011";
		Trees_din <= x"000dd210";
		wait for Clk_period;
		Addr <=  "00000111011100";
		Trees_din <= x"05fb6608";
		wait for Clk_period;
		Addr <=  "00000111011101";
		Trees_din <= x"12028704";
		wait for Clk_period;
		Addr <=  "00000111011110";
		Trees_din <= x"00d807fd";
		wait for Clk_period;
		Addr <=  "00000111011111";
		Trees_din <= x"009b07fd";
		wait for Clk_period;
		Addr <=  "00000111100000";
		Trees_din <= x"0204f604";
		wait for Clk_period;
		Addr <=  "00000111100001";
		Trees_din <= x"009007fd";
		wait for Clk_period;
		Addr <=  "00000111100010";
		Trees_din <= x"ff5c07fd";
		wait for Clk_period;
		Addr <=  "00000111100011";
		Trees_din <= x"04fd2008";
		wait for Clk_period;
		Addr <=  "00000111100100";
		Trees_din <= x"15007804";
		wait for Clk_period;
		Addr <=  "00000111100101";
		Trees_din <= x"ff7807fd";
		wait for Clk_period;
		Addr <=  "00000111100110";
		Trees_din <= x"009e07fd";
		wait for Clk_period;
		Addr <=  "00000111100111";
		Trees_din <= x"02ff4204";
		wait for Clk_period;
		Addr <=  "00000111101000";
		Trees_din <= x"00e207fd";
		wait for Clk_period;
		Addr <=  "00000111101001";
		Trees_din <= x"ff3307fd";
		wait for Clk_period;
		Addr <=  "00000111101010";
		Trees_din <= x"0112d618";
		wait for Clk_period;
		Addr <=  "00000111101011";
		Trees_din <= x"03f7f010";
		wait for Clk_period;
		Addr <=  "00000111101100";
		Trees_din <= x"1f000208";
		wait for Clk_period;
		Addr <=  "00000111101101";
		Trees_din <= x"0a079004";
		wait for Clk_period;
		Addr <=  "00000111101110";
		Trees_din <= x"ff6907fd";
		wait for Clk_period;
		Addr <=  "00000111101111";
		Trees_din <= x"003e07fd";
		wait for Clk_period;
		Addr <=  "00000111110000";
		Trees_din <= x"09005704";
		wait for Clk_period;
		Addr <=  "00000111110001";
		Trees_din <= x"ff8407fd";
		wait for Clk_period;
		Addr <=  "00000111110010";
		Trees_din <= x"00d907fd";
		wait for Clk_period;
		Addr <=  "00000111110011";
		Trees_din <= x"07005604";
		wait for Clk_period;
		Addr <=  "00000111110100";
		Trees_din <= x"00dc07fd";
		wait for Clk_period;
		Addr <=  "00000111110101";
		Trees_din <= x"ff9907fd";
		wait for Clk_period;
		Addr <=  "00000111110110";
		Trees_din <= x"0801ca08";
		wait for Clk_period;
		Addr <=  "00000111110111";
		Trees_din <= x"02016004";
		wait for Clk_period;
		Addr <=  "00000111111000";
		Trees_din <= x"003807fd";
		wait for Clk_period;
		Addr <=  "00000111111001";
		Trees_din <= x"ff7107fd";
		wait for Clk_period;
		Addr <=  "00000111111010";
		Trees_din <= x"13fe4408";
		wait for Clk_period;
		Addr <=  "00000111111011";
		Trees_din <= x"0c010104";
		wait for Clk_period;
		Addr <=  "00000111111100";
		Trees_din <= x"fff107fd";
		wait for Clk_period;
		Addr <=  "00000111111101";
		Trees_din <= x"012407fd";
		wait for Clk_period;
		Addr <=  "00000111111110";
		Trees_din <= x"ff9707fd";
		wait for Clk_period;
		Addr <=  "00000111111111";
		Trees_din <= x"01084154";
		wait for Clk_period;
		Addr <=  "00001000000000";
		Trees_din <= x"000e0e30";
		wait for Clk_period;
		Addr <=  "00001000000001";
		Trees_din <= x"01017518";
		wait for Clk_period;
		Addr <=  "00001000000010";
		Trees_din <= x"0f03e60c";
		wait for Clk_period;
		Addr <=  "00001000000011";
		Trees_din <= x"07005e04";
		wait for Clk_period;
		Addr <=  "00001000000100";
		Trees_din <= x"ff630951";
		wait for Clk_period;
		Addr <=  "00001000000101";
		Trees_din <= x"02ff0f04";
		wait for Clk_period;
		Addr <=  "00001000000110";
		Trees_din <= x"ffa90951";
		wait for Clk_period;
		Addr <=  "00001000000111";
		Trees_din <= x"00480951";
		wait for Clk_period;
		Addr <=  "00001000001000";
		Trees_din <= x"01fe5b04";
		wait for Clk_period;
		Addr <=  "00001000001001";
		Trees_din <= x"ff7a0951";
		wait for Clk_period;
		Addr <=  "00001000001010";
		Trees_din <= x"11012204";
		wait for Clk_period;
		Addr <=  "00001000001011";
		Trees_din <= x"01160951";
		wait for Clk_period;
		Addr <=  "00001000001100";
		Trees_din <= x"ff9b0951";
		wait for Clk_period;
		Addr <=  "00001000001101";
		Trees_din <= x"07005e10";
		wait for Clk_period;
		Addr <=  "00001000001110";
		Trees_din <= x"020c6008";
		wait for Clk_period;
		Addr <=  "00001000001111";
		Trees_din <= x"04fbba04";
		wait for Clk_period;
		Addr <=  "00001000010000";
		Trees_din <= x"006b0951";
		wait for Clk_period;
		Addr <=  "00001000010001";
		Trees_din <= x"ffed0951";
		wait for Clk_period;
		Addr <=  "00001000010010";
		Trees_din <= x"0f000104";
		wait for Clk_period;
		Addr <=  "00001000010011";
		Trees_din <= x"00400951";
		wait for Clk_period;
		Addr <=  "00001000010100";
		Trees_din <= x"ff670951";
		wait for Clk_period;
		Addr <=  "00001000010101";
		Trees_din <= x"08004e04";
		wait for Clk_period;
		Addr <=  "00001000010110";
		Trees_din <= x"018b0951";
		wait for Clk_period;
		Addr <=  "00001000010111";
		Trees_din <= x"004a0951";
		wait for Clk_period;
		Addr <=  "00001000011000";
		Trees_din <= x"0014ad18";
		wait for Clk_period;
		Addr <=  "00001000011001";
		Trees_din <= x"1600aa0c";
		wait for Clk_period;
		Addr <=  "00001000011010";
		Trees_din <= x"0105aa04";
		wait for Clk_period;
		Addr <=  "00001000011011";
		Trees_din <= x"ff6f0951";
		wait for Clk_period;
		Addr <=  "00001000011100";
		Trees_din <= x"0afc5304";
		wait for Clk_period;
		Addr <=  "00001000011101";
		Trees_din <= x"017c0951";
		wait for Clk_period;
		Addr <=  "00001000011110";
		Trees_din <= x"ff900951";
		wait for Clk_period;
		Addr <=  "00001000011111";
		Trees_din <= x"0f02af04";
		wait for Clk_period;
		Addr <=  "00001000100000";
		Trees_din <= x"ff620951";
		wait for Clk_period;
		Addr <=  "00001000100001";
		Trees_din <= x"07005804";
		wait for Clk_period;
		Addr <=  "00001000100010";
		Trees_din <= x"ff950951";
		wait for Clk_period;
		Addr <=  "00001000100011";
		Trees_din <= x"00490951";
		wait for Clk_period;
		Addr <=  "00001000100100";
		Trees_din <= x"0d000008";
		wait for Clk_period;
		Addr <=  "00001000100101";
		Trees_din <= x"1c003204";
		wait for Clk_period;
		Addr <=  "00001000100110";
		Trees_din <= x"00470951";
		wait for Clk_period;
		Addr <=  "00001000100111";
		Trees_din <= x"ff850951";
		wait for Clk_period;
		Addr <=  "00001000101000";
		Trees_din <= x"ff620951";
		wait for Clk_period;
		Addr <=  "00001000101001";
		Trees_din <= x"0016763c";
		wait for Clk_period;
		Addr <=  "00001000101010";
		Trees_din <= x"0111ec20";
		wait for Clk_period;
		Addr <=  "00001000101011";
		Trees_din <= x"0007fa10";
		wait for Clk_period;
		Addr <=  "00001000101100";
		Trees_din <= x"00fcaf08";
		wait for Clk_period;
		Addr <=  "00001000101101";
		Trees_din <= x"04fd2004";
		wait for Clk_period;
		Addr <=  "00001000101110";
		Trees_din <= x"007e0951";
		wait for Clk_period;
		Addr <=  "00001000101111";
		Trees_din <= x"ff8e0951";
		wait for Clk_period;
		Addr <=  "00001000110000";
		Trees_din <= x"1603df04";
		wait for Clk_period;
		Addr <=  "00001000110001";
		Trees_din <= x"00a60951";
		wait for Clk_period;
		Addr <=  "00001000110010";
		Trees_din <= x"00240951";
		wait for Clk_period;
		Addr <=  "00001000110011";
		Trees_din <= x"0c03c808";
		wait for Clk_period;
		Addr <=  "00001000110100";
		Trees_din <= x"1703f804";
		wait for Clk_period;
		Addr <=  "00001000110101";
		Trees_din <= x"00280951";
		wait for Clk_period;
		Addr <=  "00001000110110";
		Trees_din <= x"010f0951";
		wait for Clk_period;
		Addr <=  "00001000110111";
		Trees_din <= x"0b050104";
		wait for Clk_period;
		Addr <=  "00001000111000";
		Trees_din <= x"01150951";
		wait for Clk_period;
		Addr <=  "00001000111001";
		Trees_din <= x"ff930951";
		wait for Clk_period;
		Addr <=  "00001000111010";
		Trees_din <= x"02080c0c";
		wait for Clk_period;
		Addr <=  "00001000111011";
		Trees_din <= x"15007104";
		wait for Clk_period;
		Addr <=  "00001000111100";
		Trees_din <= x"ffdb0951";
		wait for Clk_period;
		Addr <=  "00001000111101";
		Trees_din <= x"000d6304";
		wait for Clk_period;
		Addr <=  "00001000111110";
		Trees_din <= x"00c10951";
		wait for Clk_period;
		Addr <=  "00001000111111";
		Trees_din <= x"00910951";
		wait for Clk_period;
		Addr <=  "00001001000000";
		Trees_din <= x"04f9df08";
		wait for Clk_period;
		Addr <=  "00001001000001";
		Trees_din <= x"12021004";
		wait for Clk_period;
		Addr <=  "00001001000010";
		Trees_din <= x"00b00951";
		wait for Clk_period;
		Addr <=  "00001001000011";
		Trees_din <= x"00140951";
		wait for Clk_period;
		Addr <=  "00001001000100";
		Trees_din <= x"04fd7904";
		wait for Clk_period;
		Addr <=  "00001001000101";
		Trees_din <= x"ff6a0951";
		wait for Clk_period;
		Addr <=  "00001001000110";
		Trees_din <= x"008f0951";
		wait for Clk_period;
		Addr <=  "00001001000111";
		Trees_din <= x"010e310c";
		wait for Clk_period;
		Addr <=  "00001001001000";
		Trees_din <= x"0c03e908";
		wait for Clk_period;
		Addr <=  "00001001001001";
		Trees_din <= x"1f000c04";
		wait for Clk_period;
		Addr <=  "00001001001010";
		Trees_din <= x"ff630951";
		wait for Clk_period;
		Addr <=  "00001001001011";
		Trees_din <= x"001b0951";
		wait for Clk_period;
		Addr <=  "00001001001100";
		Trees_din <= x"00260951";
		wait for Clk_period;
		Addr <=  "00001001001101";
		Trees_din <= x"001df30c";
		wait for Clk_period;
		Addr <=  "00001001001110";
		Trees_din <= x"17000004";
		wait for Clk_period;
		Addr <=  "00001001001111";
		Trees_din <= x"ff7b0951";
		wait for Clk_period;
		Addr <=  "00001001010000";
		Trees_din <= x"1d003e04";
		wait for Clk_period;
		Addr <=  "00001001010001";
		Trees_din <= x"ffb70951";
		wait for Clk_period;
		Addr <=  "00001001010010";
		Trees_din <= x"009c0951";
		wait for Clk_period;
		Addr <=  "00001001010011";
		Trees_din <= x"ff700951";
		wait for Clk_period;
		Addr <=  "00001001010100";
		Trees_din <= x"0108415c";
		wait for Clk_period;
		Addr <=  "00001001010101";
		Trees_din <= x"000e0e30";
		wait for Clk_period;
		Addr <=  "00001001010110";
		Trees_din <= x"01017514";
		wait for Clk_period;
		Addr <=  "00001001010111";
		Trees_din <= x"0f03e608";
		wait for Clk_period;
		Addr <=  "00001001011000";
		Trees_din <= x"07005e04";
		wait for Clk_period;
		Addr <=  "00001001011001";
		Trees_din <= x"ff660ab5";
		wait for Clk_period;
		Addr <=  "00001001011010";
		Trees_din <= x"fffe0ab5";
		wait for Clk_period;
		Addr <=  "00001001011011";
		Trees_din <= x"16001c04";
		wait for Clk_period;
		Addr <=  "00001001011100";
		Trees_din <= x"ff7f0ab5";
		wait for Clk_period;
		Addr <=  "00001001011101";
		Trees_din <= x"05fb2b04";
		wait for Clk_period;
		Addr <=  "00001001011110";
		Trees_din <= x"ffa20ab5";
		wait for Clk_period;
		Addr <=  "00001001011111";
		Trees_din <= x"00e90ab5";
		wait for Clk_period;
		Addr <=  "00001001100000";
		Trees_din <= x"07005d10";
		wait for Clk_period;
		Addr <=  "00001001100001";
		Trees_din <= x"020c6008";
		wait for Clk_period;
		Addr <=  "00001001100010";
		Trees_din <= x"1a00e204";
		wait for Clk_period;
		Addr <=  "00001001100011";
		Trees_din <= x"ffe70ab5";
		wait for Clk_period;
		Addr <=  "00001001100100";
		Trees_din <= x"004a0ab5";
		wait for Clk_period;
		Addr <=  "00001001100101";
		Trees_din <= x"0f000104";
		wait for Clk_period;
		Addr <=  "00001001100110";
		Trees_din <= x"00430ab5";
		wait for Clk_period;
		Addr <=  "00001001100111";
		Trees_din <= x"ff6b0ab5";
		wait for Clk_period;
		Addr <=  "00001001101000";
		Trees_din <= x"1b004408";
		wait for Clk_period;
		Addr <=  "00001001101001";
		Trees_din <= x"17036004";
		wait for Clk_period;
		Addr <=  "00001001101010";
		Trees_din <= x"ff920ab5";
		wait for Clk_period;
		Addr <=  "00001001101011";
		Trees_din <= x"00a70ab5";
		wait for Clk_period;
		Addr <=  "00001001101100";
		Trees_din <= x"014a0ab5";
		wait for Clk_period;
		Addr <=  "00001001101101";
		Trees_din <= x"03f87814";
		wait for Clk_period;
		Addr <=  "00001001101110";
		Trees_din <= x"0d000008";
		wait for Clk_period;
		Addr <=  "00001001101111";
		Trees_din <= x"19009b04";
		wait for Clk_period;
		Addr <=  "00001001110000";
		Trees_din <= x"ff900ab5";
		wait for Clk_period;
		Addr <=  "00001001110001";
		Trees_din <= x"00460ab5";
		wait for Clk_period;
		Addr <=  "00001001110010";
		Trees_din <= x"21000004";
		wait for Clk_period;
		Addr <=  "00001001110011";
		Trees_din <= x"ff630ab5";
		wait for Clk_period;
		Addr <=  "00001001110100";
		Trees_din <= x"1d004904";
		wait for Clk_period;
		Addr <=  "00001001110101";
		Trees_din <= x"ff7a0ab5";
		wait for Clk_period;
		Addr <=  "00001001110110";
		Trees_din <= x"00490ab5";
		wait for Clk_period;
		Addr <=  "00001001110111";
		Trees_din <= x"1600aa0c";
		wait for Clk_period;
		Addr <=  "00001001111000";
		Trees_din <= x"0105aa04";
		wait for Clk_period;
		Addr <=  "00001001111001";
		Trees_din <= x"ff740ab5";
		wait for Clk_period;
		Addr <=  "00001001111010";
		Trees_din <= x"18004204";
		wait for Clk_period;
		Addr <=  "00001001111011";
		Trees_din <= x"01800ab5";
		wait for Clk_period;
		Addr <=  "00001001111100";
		Trees_din <= x"ff9d0ab5";
		wait for Clk_period;
		Addr <=  "00001001111101";
		Trees_din <= x"0f02af04";
		wait for Clk_period;
		Addr <=  "00001001111110";
		Trees_din <= x"ff650ab5";
		wait for Clk_period;
		Addr <=  "00001001111111";
		Trees_din <= x"1b003b04";
		wait for Clk_period;
		Addr <=  "00001010000000";
		Trees_din <= x"ff960ab5";
		wait for Clk_period;
		Addr <=  "00001010000001";
		Trees_din <= x"00480ab5";
		wait for Clk_period;
		Addr <=  "00001010000010";
		Trees_din <= x"00167638";
		wait for Clk_period;
		Addr <=  "00001010000011";
		Trees_din <= x"0113e920";
		wait for Clk_period;
		Addr <=  "00001010000100";
		Trees_din <= x"0007fa10";
		wait for Clk_period;
		Addr <=  "00001010000101";
		Trees_din <= x"010a4208";
		wait for Clk_period;
		Addr <=  "00001010000110";
		Trees_din <= x"1d004e04";
		wait for Clk_period;
		Addr <=  "00001010000111";
		Trees_din <= x"fffe0ab5";
		wait for Clk_period;
		Addr <=  "00001010001000";
		Trees_din <= x"00c30ab5";
		wait for Clk_period;
		Addr <=  "00001010001001";
		Trees_din <= x"14001d04";
		wait for Clk_period;
		Addr <=  "00001010001010";
		Trees_din <= x"ffc00ab5";
		wait for Clk_period;
		Addr <=  "00001010001011";
		Trees_din <= x"00900ab5";
		wait for Clk_period;
		Addr <=  "00001010001100";
		Trees_din <= x"0afccc08";
		wait for Clk_period;
		Addr <=  "00001010001101";
		Trees_din <= x"010fd304";
		wait for Clk_period;
		Addr <=  "00001010001110";
		Trees_din <= x"00360ab5";
		wait for Clk_period;
		Addr <=  "00001010001111";
		Trees_din <= x"00950ab5";
		wait for Clk_period;
		Addr <=  "00001010010000";
		Trees_din <= x"16000504";
		wait for Clk_period;
		Addr <=  "00001010010001";
		Trees_din <= x"ff6d0ab5";
		wait for Clk_period;
		Addr <=  "00001010010010";
		Trees_din <= x"00210ab5";
		wait for Clk_period;
		Addr <=  "00001010010011";
		Trees_din <= x"0013bd0c";
		wait for Clk_period;
		Addr <=  "00001010010100";
		Trees_din <= x"22000008";
		wait for Clk_period;
		Addr <=  "00001010010101";
		Trees_din <= x"0ef98004";
		wait for Clk_period;
		Addr <=  "00001010010110";
		Trees_din <= x"003e0ab5";
		wait for Clk_period;
		Addr <=  "00001010010111";
		Trees_din <= x"00bc0ab5";
		wait for Clk_period;
		Addr <=  "00001010011000";
		Trees_din <= x"ffec0ab5";
		wait for Clk_period;
		Addr <=  "00001010011001";
		Trees_din <= x"07005504";
		wait for Clk_period;
		Addr <=  "00001010011010";
		Trees_din <= x"ffa10ab5";
		wait for Clk_period;
		Addr <=  "00001010011011";
		Trees_din <= x"1201b904";
		wait for Clk_period;
		Addr <=  "00001010011100";
		Trees_din <= x"00b70ab5";
		wait for Clk_period;
		Addr <=  "00001010011101";
		Trees_din <= x"ffe90ab5";
		wait for Clk_period;
		Addr <=  "00001010011110";
		Trees_din <= x"010e310c";
		wait for Clk_period;
		Addr <=  "00001010011111";
		Trees_din <= x"0c03e908";
		wait for Clk_period;
		Addr <=  "00001010100000";
		Trees_din <= x"1f000c04";
		wait for Clk_period;
		Addr <=  "00001010100001";
		Trees_din <= x"ff660ab5";
		wait for Clk_period;
		Addr <=  "00001010100010";
		Trees_din <= x"00260ab5";
		wait for Clk_period;
		Addr <=  "00001010100011";
		Trees_din <= x"002a0ab5";
		wait for Clk_period;
		Addr <=  "00001010100100";
		Trees_din <= x"001df310";
		wait for Clk_period;
		Addr <=  "00001010100101";
		Trees_din <= x"07005508";
		wait for Clk_period;
		Addr <=  "00001010100110";
		Trees_din <= x"06f50204";
		wait for Clk_period;
		Addr <=  "00001010100111";
		Trees_din <= x"00e00ab5";
		wait for Clk_period;
		Addr <=  "00001010101000";
		Trees_din <= x"ff9c0ab5";
		wait for Clk_period;
		Addr <=  "00001010101001";
		Trees_din <= x"0d031e04";
		wait for Clk_period;
		Addr <=  "00001010101010";
		Trees_din <= x"ff860ab5";
		wait for Clk_period;
		Addr <=  "00001010101011";
		Trees_din <= x"008e0ab5";
		wait for Clk_period;
		Addr <=  "00001010101100";
		Trees_din <= x"ff760ab5";
		wait for Clk_period;
		Addr <=  "00001010101101";
		Trees_din <= x"0105bc4c";
		wait for Clk_period;
		Addr <=  "00001010101110";
		Trees_din <= x"03fc9714";
		wait for Clk_period;
		Addr <=  "00001010101111";
		Trees_din <= x"16040010";
		wait for Clk_period;
		Addr <=  "00001010110000";
		Trees_din <= x"0105aa0c";
		wait for Clk_period;
		Addr <=  "00001010110001";
		Trees_din <= x"0d000008";
		wait for Clk_period;
		Addr <=  "00001010110010";
		Trees_din <= x"0a027804";
		wait for Clk_period;
		Addr <=  "00001010110011";
		Trees_din <= x"00490c19";
		wait for Clk_period;
		Addr <=  "00001010110100";
		Trees_din <= x"ff9c0c19";
		wait for Clk_period;
		Addr <=  "00001010110101";
		Trees_din <= x"ff640c19";
		wait for Clk_period;
		Addr <=  "00001010110110";
		Trees_din <= x"002e0c19";
		wait for Clk_period;
		Addr <=  "00001010110111";
		Trees_din <= x"003b0c19";
		wait for Clk_period;
		Addr <=  "00001010111000";
		Trees_din <= x"01017518";
		wait for Clk_period;
		Addr <=  "00001010111001";
		Trees_din <= x"0f03e60c";
		wait for Clk_period;
		Addr <=  "00001010111010";
		Trees_din <= x"07005e08";
		wait for Clk_period;
		Addr <=  "00001010111011";
		Trees_din <= x"0af83804";
		wait for Clk_period;
		Addr <=  "00001010111100";
		Trees_din <= x"ffa00c19";
		wait for Clk_period;
		Addr <=  "00001010111101";
		Trees_din <= x"ff640c19";
		wait for Clk_period;
		Addr <=  "00001010111110";
		Trees_din <= x"00190c19";
		wait for Clk_period;
		Addr <=  "00001010111111";
		Trees_din <= x"01fe4904";
		wait for Clk_period;
		Addr <=  "00001011000000";
		Trees_din <= x"ff860c19";
		wait for Clk_period;
		Addr <=  "00001011000001";
		Trees_din <= x"16001804";
		wait for Clk_period;
		Addr <=  "00001011000010";
		Trees_din <= x"ffae0c19";
		wait for Clk_period;
		Addr <=  "00001011000011";
		Trees_din <= x"00d30c19";
		wait for Clk_period;
		Addr <=  "00001011000100";
		Trees_din <= x"0d02c810";
		wait for Clk_period;
		Addr <=  "00001011000101";
		Trees_din <= x"1d003708";
		wait for Clk_period;
		Addr <=  "00001011000110";
		Trees_din <= x"1900b404";
		wait for Clk_period;
		Addr <=  "00001011000111";
		Trees_din <= x"00fd0c19";
		wait for Clk_period;
		Addr <=  "00001011001000";
		Trees_din <= x"ff870c19";
		wait for Clk_period;
		Addr <=  "00001011001001";
		Trees_din <= x"08000504";
		wait for Clk_period;
		Addr <=  "00001011001010";
		Trees_din <= x"00990c19";
		wait for Clk_period;
		Addr <=  "00001011001011";
		Trees_din <= x"ff970c19";
		wait for Clk_period;
		Addr <=  "00001011001100";
		Trees_din <= x"04fb2808";
		wait for Clk_period;
		Addr <=  "00001011001101";
		Trees_din <= x"1b003704";
		wait for Clk_period;
		Addr <=  "00001011001110";
		Trees_din <= x"ff9c0c19";
		wait for Clk_period;
		Addr <=  "00001011001111";
		Trees_din <= x"023b0c19";
		wait for Clk_period;
		Addr <=  "00001011010000";
		Trees_din <= x"03fe8b04";
		wait for Clk_period;
		Addr <=  "00001011010001";
		Trees_din <= x"012d0c19";
		wait for Clk_period;
		Addr <=  "00001011010010";
		Trees_din <= x"ffbc0c19";
		wait for Clk_period;
		Addr <=  "00001011010011";
		Trees_din <= x"00173a3c";
		wait for Clk_period;
		Addr <=  "00001011010100";
		Trees_din <= x"010d4f20";
		wait for Clk_period;
		Addr <=  "00001011010101";
		Trees_din <= x"03f6f410";
		wait for Clk_period;
		Addr <=  "00001011010110";
		Trees_din <= x"10fa8508";
		wait for Clk_period;
		Addr <=  "00001011010111";
		Trees_din <= x"04f99004";
		wait for Clk_period;
		Addr <=  "00001011011000";
		Trees_din <= x"ff8c0c19";
		wait for Clk_period;
		Addr <=  "00001011011001";
		Trees_din <= x"00d40c19";
		wait for Clk_period;
		Addr <=  "00001011011010";
		Trees_din <= x"04f81504";
		wait for Clk_period;
		Addr <=  "00001011011011";
		Trees_din <= x"ffbe0c19";
		wait for Clk_period;
		Addr <=  "00001011011100";
		Trees_din <= x"ff5b0c19";
		wait for Clk_period;
		Addr <=  "00001011011101";
		Trees_din <= x"010d2808";
		wait for Clk_period;
		Addr <=  "00001011011110";
		Trees_din <= x"010cb404";
		wait for Clk_period;
		Addr <=  "00001011011111";
		Trees_din <= x"00270c19";
		wait for Clk_period;
		Addr <=  "00001011100000";
		Trees_din <= x"009c0c19";
		wait for Clk_period;
		Addr <=  "00001011100001";
		Trees_din <= x"14031004";
		wait for Clk_period;
		Addr <=  "00001011100010";
		Trees_din <= x"ff360c19";
		wait for Clk_period;
		Addr <=  "00001011100011";
		Trees_din <= x"00050c19";
		wait for Clk_period;
		Addr <=  "00001011100100";
		Trees_din <= x"01159310";
		wait for Clk_period;
		Addr <=  "00001011100101";
		Trees_din <= x"03f9d608";
		wait for Clk_period;
		Addr <=  "00001011100110";
		Trees_din <= x"06f66004";
		wait for Clk_period;
		Addr <=  "00001011100111";
		Trees_din <= x"00250c19";
		wait for Clk_period;
		Addr <=  "00001011101000";
		Trees_din <= x"00750c19";
		wait for Clk_period;
		Addr <=  "00001011101001";
		Trees_din <= x"05f98f04";
		wait for Clk_period;
		Addr <=  "00001011101010";
		Trees_din <= x"00590c19";
		wait for Clk_period;
		Addr <=  "00001011101011";
		Trees_din <= x"00b40c19";
		wait for Clk_period;
		Addr <=  "00001011101100";
		Trees_din <= x"21000008";
		wait for Clk_period;
		Addr <=  "00001011101101";
		Trees_din <= x"020a1904";
		wait for Clk_period;
		Addr <=  "00001011101110";
		Trees_din <= x"00ae0c19";
		wait for Clk_period;
		Addr <=  "00001011101111";
		Trees_din <= x"00270c19";
		wait for Clk_period;
		Addr <=  "00001011110000";
		Trees_din <= x"000c0c19";
		wait for Clk_period;
		Addr <=  "00001011110001";
		Trees_din <= x"0112d618";
		wait for Clk_period;
		Addr <=  "00001011110010";
		Trees_din <= x"07004808";
		wait for Clk_period;
		Addr <=  "00001011110011";
		Trees_din <= x"1d004804";
		wait for Clk_period;
		Addr <=  "00001011110100";
		Trees_din <= x"ffa40c19";
		wait for Clk_period;
		Addr <=  "00001011110101";
		Trees_din <= x"00d60c19";
		wait for Clk_period;
		Addr <=  "00001011110110";
		Trees_din <= x"11043808";
		wait for Clk_period;
		Addr <=  "00001011110111";
		Trees_din <= x"1f000c04";
		wait for Clk_period;
		Addr <=  "00001011111000";
		Trees_din <= x"ff6c0c19";
		wait for Clk_period;
		Addr <=  "00001011111001";
		Trees_din <= x"00120c19";
		wait for Clk_period;
		Addr <=  "00001011111010";
		Trees_din <= x"11045604";
		wait for Clk_period;
		Addr <=  "00001011111011";
		Trees_din <= x"00960c19";
		wait for Clk_period;
		Addr <=  "00001011111100";
		Trees_din <= x"ff820c19";
		wait for Clk_period;
		Addr <=  "00001011111101";
		Trees_din <= x"0801ca08";
		wait for Clk_period;
		Addr <=  "00001011111110";
		Trees_din <= x"1103d604";
		wait for Clk_period;
		Addr <=  "00001011111111";
		Trees_din <= x"ff820c19";
		wait for Clk_period;
		Addr <=  "00001100000000";
		Trees_din <= x"00270c19";
		wait for Clk_period;
		Addr <=  "00001100000001";
		Trees_din <= x"0c010104";
		wait for Clk_period;
		Addr <=  "00001100000010";
		Trees_din <= x"fff10c19";
		wait for Clk_period;
		Addr <=  "00001100000011";
		Trees_din <= x"14018a04";
		wait for Clk_period;
		Addr <=  "00001100000100";
		Trees_din <= x"00dd0c19";
		wait for Clk_period;
		Addr <=  "00001100000101";
		Trees_din <= x"00140c19";
		wait for Clk_period;
		Addr <=  "00001100000110";
		Trees_din <= x"0105bc48";
		wait for Clk_period;
		Addr <=  "00001100000111";
		Trees_din <= x"03fc9714";
		wait for Clk_period;
		Addr <=  "00001100001000";
		Trees_din <= x"0105aa10";
		wait for Clk_period;
		Addr <=  "00001100001001";
		Trees_din <= x"14000b04";
		wait for Clk_period;
		Addr <=  "00001100001010";
		Trees_din <= x"00230d5d";
		wait for Clk_period;
		Addr <=  "00001100001011";
		Trees_din <= x"0d000008";
		wait for Clk_period;
		Addr <=  "00001100001100";
		Trees_din <= x"09005404";
		wait for Clk_period;
		Addr <=  "00001100001101";
		Trees_din <= x"004a0d5d";
		wait for Clk_period;
		Addr <=  "00001100001110";
		Trees_din <= x"ffa60d5d";
		wait for Clk_period;
		Addr <=  "00001100001111";
		Trees_din <= x"ff650d5d";
		wait for Clk_period;
		Addr <=  "00001100010000";
		Trees_din <= x"00340d5d";
		wait for Clk_period;
		Addr <=  "00001100010001";
		Trees_din <= x"01017518";
		wait for Clk_period;
		Addr <=  "00001100010010";
		Trees_din <= x"0f03e60c";
		wait for Clk_period;
		Addr <=  "00001100010011";
		Trees_din <= x"07005e08";
		wait for Clk_period;
		Addr <=  "00001100010100";
		Trees_din <= x"05ff4a04";
		wait for Clk_period;
		Addr <=  "00001100010101";
		Trees_din <= x"ff660d5d";
		wait for Clk_period;
		Addr <=  "00001100010110";
		Trees_din <= x"ffa90d5d";
		wait for Clk_period;
		Addr <=  "00001100010111";
		Trees_din <= x"00200d5d";
		wait for Clk_period;
		Addr <=  "00001100011000";
		Trees_din <= x"01fe4904";
		wait for Clk_period;
		Addr <=  "00001100011001";
		Trees_din <= x"ff8c0d5d";
		wait for Clk_period;
		Addr <=  "00001100011010";
		Trees_din <= x"0efee804";
		wait for Clk_period;
		Addr <=  "00001100011011";
		Trees_din <= x"ffab0d5d";
		wait for Clk_period;
		Addr <=  "00001100011100";
		Trees_din <= x"00bc0d5d";
		wait for Clk_period;
		Addr <=  "00001100011101";
		Trees_din <= x"0c036410";
		wait for Clk_period;
		Addr <=  "00001100011110";
		Trees_din <= x"19009e08";
		wait for Clk_period;
		Addr <=  "00001100011111";
		Trees_din <= x"06fb2904";
		wait for Clk_period;
		Addr <=  "00001100100000";
		Trees_din <= x"ff830d5d";
		wait for Clk_period;
		Addr <=  "00001100100001";
		Trees_din <= x"007b0d5d";
		wait for Clk_period;
		Addr <=  "00001100100010";
		Trees_din <= x"19009f04";
		wait for Clk_period;
		Addr <=  "00001100100011";
		Trees_din <= x"01c90d5d";
		wait for Clk_period;
		Addr <=  "00001100100100";
		Trees_din <= x"000f0d5d";
		wait for Clk_period;
		Addr <=  "00001100100101";
		Trees_din <= x"09005908";
		wait for Clk_period;
		Addr <=  "00001100100110";
		Trees_din <= x"1500ad04";
		wait for Clk_period;
		Addr <=  "00001100100111";
		Trees_din <= x"ffa40d5d";
		wait for Clk_period;
		Addr <=  "00001100101000";
		Trees_din <= x"013f0d5d";
		wait for Clk_period;
		Addr <=  "00001100101001";
		Trees_din <= x"01550d5d";
		wait for Clk_period;
		Addr <=  "00001100101010";
		Trees_din <= x"0018d040";
		wait for Clk_period;
		Addr <=  "00001100101011";
		Trees_din <= x"0113e920";
		wait for Clk_period;
		Addr <=  "00001100101100";
		Trees_din <= x"010c8d10";
		wait for Clk_period;
		Addr <=  "00001100101101";
		Trees_din <= x"03f6f408";
		wait for Clk_period;
		Addr <=  "00001100101110";
		Trees_din <= x"09005c04";
		wait for Clk_period;
		Addr <=  "00001100101111";
		Trees_din <= x"ff670d5d";
		wait for Clk_period;
		Addr <=  "00001100110000";
		Trees_din <= x"00880d5d";
		wait for Clk_period;
		Addr <=  "00001100110001";
		Trees_din <= x"11032704";
		wait for Clk_period;
		Addr <=  "00001100110010";
		Trees_din <= x"002f0d5d";
		wait for Clk_period;
		Addr <=  "00001100110011";
		Trees_din <= x"ffdc0d5d";
		wait for Clk_period;
		Addr <=  "00001100110100";
		Trees_din <= x"0a000e08";
		wait for Clk_period;
		Addr <=  "00001100110101";
		Trees_din <= x"0802ad04";
		wait for Clk_period;
		Addr <=  "00001100110110";
		Trees_din <= x"00500d5d";
		wait for Clk_period;
		Addr <=  "00001100110111";
		Trees_din <= x"00de0d5d";
		wait for Clk_period;
		Addr <=  "00001100111000";
		Trees_din <= x"0003aa04";
		wait for Clk_period;
		Addr <=  "00001100111001";
		Trees_din <= x"008b0d5d";
		wait for Clk_period;
		Addr <=  "00001100111010";
		Trees_din <= x"00100d5d";
		wait for Clk_period;
		Addr <=  "00001100111011";
		Trees_din <= x"0013bd10";
		wait for Clk_period;
		Addr <=  "00001100111100";
		Trees_din <= x"0ef98008";
		wait for Clk_period;
		Addr <=  "00001100111101";
		Trees_din <= x"03f68204";
		wait for Clk_period;
		Addr <=  "00001100111110";
		Trees_din <= x"ff8a0d5d";
		wait for Clk_period;
		Addr <=  "00001100111111";
		Trees_din <= x"007c0d5d";
		wait for Clk_period;
		Addr <=  "00001101000000";
		Trees_din <= x"22000004";
		wait for Clk_period;
		Addr <=  "00001101000001";
		Trees_din <= x"00a70d5d";
		wait for Clk_period;
		Addr <=  "00001101000010";
		Trees_din <= x"ffe50d5d";
		wait for Clk_period;
		Addr <=  "00001101000011";
		Trees_din <= x"10fb3708";
		wait for Clk_period;
		Addr <=  "00001101000100";
		Trees_din <= x"09005404";
		wait for Clk_period;
		Addr <=  "00001101000101";
		Trees_din <= x"00070d5d";
		wait for Clk_period;
		Addr <=  "00001101000110";
		Trees_din <= x"ff6d0d5d";
		wait for Clk_period;
		Addr <=  "00001101000111";
		Trees_din <= x"0b028804";
		wait for Clk_period;
		Addr <=  "00001101001000";
		Trees_din <= x"00b80d5d";
		wait for Clk_period;
		Addr <=  "00001101001001";
		Trees_din <= x"00000d5d";
		wait for Clk_period;
		Addr <=  "00001101001010";
		Trees_din <= x"010ed00c";
		wait for Clk_period;
		Addr <=  "00001101001011";
		Trees_din <= x"1f000c08";
		wait for Clk_period;
		Addr <=  "00001101001100";
		Trees_din <= x"21000004";
		wait for Clk_period;
		Addr <=  "00001101001101";
		Trees_din <= x"ff690d5d";
		wait for Clk_period;
		Addr <=  "00001101001110";
		Trees_din <= x"00390d5d";
		wait for Clk_period;
		Addr <=  "00001101001111";
		Trees_din <= x"002b0d5d";
		wait for Clk_period;
		Addr <=  "00001101010000";
		Trees_din <= x"1e006a04";
		wait for Clk_period;
		Addr <=  "00001101010001";
		Trees_din <= x"ff7c0d5d";
		wait for Clk_period;
		Addr <=  "00001101010010";
		Trees_din <= x"1a00b804";
		wait for Clk_period;
		Addr <=  "00001101010011";
		Trees_din <= x"ff8c0d5d";
		wait for Clk_period;
		Addr <=  "00001101010100";
		Trees_din <= x"13fdc604";
		wait for Clk_period;
		Addr <=  "00001101010101";
		Trees_din <= x"ffe90d5d";
		wait for Clk_period;
		Addr <=  "00001101010110";
		Trees_din <= x"01000d5d";
		wait for Clk_period;
		Addr <=  "00001101010111";
		Trees_din <= x"0105bc44";
		wait for Clk_period;
		Addr <=  "00001101011000";
		Trees_din <= x"03fc9714";
		wait for Clk_period;
		Addr <=  "00001101011001";
		Trees_din <= x"0105aa10";
		wait for Clk_period;
		Addr <=  "00001101011010";
		Trees_din <= x"14000b04";
		wait for Clk_period;
		Addr <=  "00001101011011";
		Trees_din <= x"002a0e89";
		wait for Clk_period;
		Addr <=  "00001101011100";
		Trees_din <= x"0d000008";
		wait for Clk_period;
		Addr <=  "00001101011101";
		Trees_din <= x"02004a04";
		wait for Clk_period;
		Addr <=  "00001101011110";
		Trees_din <= x"004a0e89";
		wait for Clk_period;
		Addr <=  "00001101011111";
		Trees_din <= x"ffb10e89";
		wait for Clk_period;
		Addr <=  "00001101100000";
		Trees_din <= x"ff660e89";
		wait for Clk_period;
		Addr <=  "00001101100001";
		Trees_din <= x"003a0e89";
		wait for Clk_period;
		Addr <=  "00001101100010";
		Trees_din <= x"01017518";
		wait for Clk_period;
		Addr <=  "00001101100011";
		Trees_din <= x"0f03e60c";
		wait for Clk_period;
		Addr <=  "00001101100100";
		Trees_din <= x"020d0608";
		wait for Clk_period;
		Addr <=  "00001101100101";
		Trees_din <= x"0af83804";
		wait for Clk_period;
		Addr <=  "00001101100110";
		Trees_din <= x"ffb40e89";
		wait for Clk_period;
		Addr <=  "00001101100111";
		Trees_din <= x"ff670e89";
		wait for Clk_period;
		Addr <=  "00001101101000";
		Trees_din <= x"00310e89";
		wait for Clk_period;
		Addr <=  "00001101101001";
		Trees_din <= x"01fe4904";
		wait for Clk_period;
		Addr <=  "00001101101010";
		Trees_din <= x"ff920e89";
		wait for Clk_period;
		Addr <=  "00001101101011";
		Trees_din <= x"03033004";
		wait for Clk_period;
		Addr <=  "00001101101100";
		Trees_din <= x"ffe10e89";
		wait for Clk_period;
		Addr <=  "00001101101101";
		Trees_din <= x"00ac0e89";
		wait for Clk_period;
		Addr <=  "00001101101110";
		Trees_din <= x"17000008";
		wait for Clk_period;
		Addr <=  "00001101101111";
		Trees_din <= x"0802df04";
		wait for Clk_period;
		Addr <=  "00001101110000";
		Trees_din <= x"ff6b0e89";
		wait for Clk_period;
		Addr <=  "00001101110001";
		Trees_din <= x"00b20e89";
		wait for Clk_period;
		Addr <=  "00001101110010";
		Trees_din <= x"0c036408";
		wait for Clk_period;
		Addr <=  "00001101110011";
		Trees_din <= x"05fa6004";
		wait for Clk_period;
		Addr <=  "00001101110100";
		Trees_din <= x"ff830e89";
		wait for Clk_period;
		Addr <=  "00001101110101";
		Trees_din <= x"003b0e89";
		wait for Clk_period;
		Addr <=  "00001101110110";
		Trees_din <= x"1b003604";
		wait for Clk_period;
		Addr <=  "00001101110111";
		Trees_din <= x"00040e89";
		wait for Clk_period;
		Addr <=  "00001101111000";
		Trees_din <= x"010d0e89";
		wait for Clk_period;
		Addr <=  "00001101111001";
		Trees_din <= x"0018d038";
		wait for Clk_period;
		Addr <=  "00001101111010";
		Trees_din <= x"0113e918";
		wait for Clk_period;
		Addr <=  "00001101111011";
		Trees_din <= x"09005e10";
		wait for Clk_period;
		Addr <=  "00001101111100";
		Trees_din <= x"15009908";
		wait for Clk_period;
		Addr <=  "00001101111101";
		Trees_din <= x"03ff5404";
		wait for Clk_period;
		Addr <=  "00001101111110";
		Trees_din <= x"002d0e89";
		wait for Clk_period;
		Addr <=  "00001101111111";
		Trees_din <= x"00850e89";
		wait for Clk_period;
		Addr <=  "00001110000000";
		Trees_din <= x"01096904";
		wait for Clk_period;
		Addr <=  "00001110000001";
		Trees_din <= x"ffd60e89";
		wait for Clk_period;
		Addr <=  "00001110000010";
		Trees_din <= x"002c0e89";
		wait for Clk_period;
		Addr <=  "00001110000011";
		Trees_din <= x"07005604";
		wait for Clk_period;
		Addr <=  "00001110000100";
		Trees_din <= x"00000e89";
		wait for Clk_period;
		Addr <=  "00001110000101";
		Trees_din <= x"ff4e0e89";
		wait for Clk_period;
		Addr <=  "00001110000110";
		Trees_din <= x"0013bd10";
		wait for Clk_period;
		Addr <=  "00001110000111";
		Trees_din <= x"0ef98008";
		wait for Clk_period;
		Addr <=  "00001110001000";
		Trees_din <= x"03f68204";
		wait for Clk_period;
		Addr <=  "00001110001001";
		Trees_din <= x"ff8e0e89";
		wait for Clk_period;
		Addr <=  "00001110001010";
		Trees_din <= x"00730e89";
		wait for Clk_period;
		Addr <=  "00001110001011";
		Trees_din <= x"020a1904";
		wait for Clk_period;
		Addr <=  "00001110001100";
		Trees_din <= x"00a30e89";
		wait for Clk_period;
		Addr <=  "00001110001101";
		Trees_din <= x"fffe0e89";
		wait for Clk_period;
		Addr <=  "00001110001110";
		Trees_din <= x"10fb3708";
		wait for Clk_period;
		Addr <=  "00001110001111";
		Trees_din <= x"09005404";
		wait for Clk_period;
		Addr <=  "00001110010000";
		Trees_din <= x"00070e89";
		wait for Clk_period;
		Addr <=  "00001110010001";
		Trees_din <= x"ff790e89";
		wait for Clk_period;
		Addr <=  "00001110010010";
		Trees_din <= x"0b028804";
		wait for Clk_period;
		Addr <=  "00001110010011";
		Trees_din <= x"00a90e89";
		wait for Clk_period;
		Addr <=  "00001110010100";
		Trees_din <= x"00060e89";
		wait for Clk_period;
		Addr <=  "00001110010101";
		Trees_din <= x"010ed00c";
		wait for Clk_period;
		Addr <=  "00001110010110";
		Trees_din <= x"0e043e08";
		wait for Clk_period;
		Addr <=  "00001110010111";
		Trees_din <= x"1f000c04";
		wait for Clk_period;
		Addr <=  "00001110011000";
		Trees_din <= x"ff6b0e89";
		wait for Clk_period;
		Addr <=  "00001110011001";
		Trees_din <= x"00350e89";
		wait for Clk_period;
		Addr <=  "00001110011010";
		Trees_din <= x"00400e89";
		wait for Clk_period;
		Addr <=  "00001110011011";
		Trees_din <= x"1d004304";
		wait for Clk_period;
		Addr <=  "00001110011100";
		Trees_din <= x"ff820e89";
		wait for Clk_period;
		Addr <=  "00001110011101";
		Trees_din <= x"1a00b804";
		wait for Clk_period;
		Addr <=  "00001110011110";
		Trees_din <= x"ff940e89";
		wait for Clk_period;
		Addr <=  "00001110011111";
		Trees_din <= x"0201e304";
		wait for Clk_period;
		Addr <=  "00001110100000";
		Trees_din <= x"013d0e89";
		wait for Clk_period;
		Addr <=  "00001110100001";
		Trees_din <= x"00250e89";
		wait for Clk_period;
		Addr <=  "00001110100010";
		Trees_din <= x"0104a624";
		wait for Clk_period;
		Addr <=  "00001110100011";
		Trees_din <= x"03fcb70c";
		wait for Clk_period;
		Addr <=  "00001110100100";
		Trees_din <= x"14000b04";
		wait for Clk_period;
		Addr <=  "00001110100101";
		Trees_din <= x"003d0f65";
		wait for Clk_period;
		Addr <=  "00001110100110";
		Trees_din <= x"0d000004";
		wait for Clk_period;
		Addr <=  "00001110100111";
		Trees_din <= x"00150f65";
		wait for Clk_period;
		Addr <=  "00001110101000";
		Trees_din <= x"ff670f65";
		wait for Clk_period;
		Addr <=  "00001110101001";
		Trees_din <= x"01fe6a04";
		wait for Clk_period;
		Addr <=  "00001110101010";
		Trees_din <= x"ff6a0f65";
		wait for Clk_period;
		Addr <=  "00001110101011";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00001110101100";
		Trees_din <= x"ff710f65";
		wait for Clk_period;
		Addr <=  "00001110101101";
		Trees_din <= x"0401dd08";
		wait for Clk_period;
		Addr <=  "00001110101110";
		Trees_din <= x"10046104";
		wait for Clk_period;
		Addr <=  "00001110101111";
		Trees_din <= x"fffd0f65";
		wait for Clk_period;
		Addr <=  "00001110110000";
		Trees_din <= x"00a00f65";
		wait for Clk_period;
		Addr <=  "00001110110001";
		Trees_din <= x"1d003704";
		wait for Clk_period;
		Addr <=  "00001110110010";
		Trees_din <= x"005d0f65";
		wait for Clk_period;
		Addr <=  "00001110110011";
		Trees_din <= x"ffb00f65";
		wait for Clk_period;
		Addr <=  "00001110110100";
		Trees_din <= x"0018d030";
		wait for Clk_period;
		Addr <=  "00001110110101";
		Trees_din <= x"01159320";
		wait for Clk_period;
		Addr <=  "00001110110110";
		Trees_din <= x"06f63b10";
		wait for Clk_period;
		Addr <=  "00001110110111";
		Trees_din <= x"06f5dc08";
		wait for Clk_period;
		Addr <=  "00001110111000";
		Trees_din <= x"1c003204";
		wait for Clk_period;
		Addr <=  "00001110111001";
		Trees_din <= x"fff70f65";
		wait for Clk_period;
		Addr <=  "00001110111010";
		Trees_din <= x"002f0f65";
		wait for Clk_period;
		Addr <=  "00001110111011";
		Trees_din <= x"010fd304";
		wait for Clk_period;
		Addr <=  "00001110111100";
		Trees_din <= x"ff7d0f65";
		wait for Clk_period;
		Addr <=  "00001110111101";
		Trees_din <= x"001a0f65";
		wait for Clk_period;
		Addr <=  "00001110111110";
		Trees_din <= x"13016508";
		wait for Clk_period;
		Addr <=  "00001110111111";
		Trees_din <= x"0104ee04";
		wait for Clk_period;
		Addr <=  "00001111000000";
		Trees_din <= x"012f0f65";
		wait for Clk_period;
		Addr <=  "00001111000001";
		Trees_din <= x"00460f65";
		wait for Clk_period;
		Addr <=  "00001111000010";
		Trees_din <= x"010b1104";
		wait for Clk_period;
		Addr <=  "00001111000011";
		Trees_din <= x"ff8a0f65";
		wait for Clk_period;
		Addr <=  "00001111000100";
		Trees_din <= x"002e0f65";
		wait for Clk_period;
		Addr <=  "00001111000101";
		Trees_din <= x"08000104";
		wait for Clk_period;
		Addr <=  "00001111000110";
		Trees_din <= x"fff20f65";
		wait for Clk_period;
		Addr <=  "00001111000111";
		Trees_din <= x"0209bd08";
		wait for Clk_period;
		Addr <=  "00001111001000";
		Trees_din <= x"10f75604";
		wait for Clk_period;
		Addr <=  "00001111001001";
		Trees_din <= x"00340f65";
		wait for Clk_period;
		Addr <=  "00001111001010";
		Trees_din <= x"00a00f65";
		wait for Clk_period;
		Addr <=  "00001111001011";
		Trees_din <= x"00060f65";
		wait for Clk_period;
		Addr <=  "00001111001100";
		Trees_din <= x"010ed00c";
		wait for Clk_period;
		Addr <=  "00001111001101";
		Trees_din <= x"09005904";
		wait for Clk_period;
		Addr <=  "00001111001110";
		Trees_din <= x"ff6c0f65";
		wait for Clk_period;
		Addr <=  "00001111001111";
		Trees_din <= x"0f02d604";
		wait for Clk_period;
		Addr <=  "00001111010000";
		Trees_din <= x"ff8b0f65";
		wait for Clk_period;
		Addr <=  "00001111010001";
		Trees_din <= x"00d00f65";
		wait for Clk_period;
		Addr <=  "00001111010010";
		Trees_din <= x"1d004304";
		wait for Clk_period;
		Addr <=  "00001111010011";
		Trees_din <= x"ff880f65";
		wait for Clk_period;
		Addr <=  "00001111010100";
		Trees_din <= x"1a00b804";
		wait for Clk_period;
		Addr <=  "00001111010101";
		Trees_din <= x"ff9b0f65";
		wait for Clk_period;
		Addr <=  "00001111010110";
		Trees_din <= x"0201e304";
		wait for Clk_period;
		Addr <=  "00001111010111";
		Trees_din <= x"01140f65";
		wait for Clk_period;
		Addr <=  "00001111011000";
		Trees_din <= x"00240f65";
		wait for Clk_period;
		Addr <=  "00001111011001";
		Trees_din <= x"0101751c";
		wait for Clk_period;
		Addr <=  "00001111011010";
		Trees_din <= x"1303b418";
		wait for Clk_period;
		Addr <=  "00001111011011";
		Trees_din <= x"07005e14";
		wait for Clk_period;
		Addr <=  "00001111011100";
		Trees_din <= x"09005e10";
		wait for Clk_period;
		Addr <=  "00001111011101";
		Trees_din <= x"06f35808";
		wait for Clk_period;
		Addr <=  "00001111011110";
		Trees_din <= x"13016804";
		wait for Clk_period;
		Addr <=  "00001111011111";
		Trees_din <= x"ff881041";
		wait for Clk_period;
		Addr <=  "00001111100000";
		Trees_din <= x"00301041";
		wait for Clk_period;
		Addr <=  "00001111100001";
		Trees_din <= x"0af83804";
		wait for Clk_period;
		Addr <=  "00001111100010";
		Trees_din <= x"ffa21041";
		wait for Clk_period;
		Addr <=  "00001111100011";
		Trees_din <= x"ff671041";
		wait for Clk_period;
		Addr <=  "00001111100100";
		Trees_din <= x"00141041";
		wait for Clk_period;
		Addr <=  "00001111100101";
		Trees_din <= x"fffd1041";
		wait for Clk_period;
		Addr <=  "00001111100110";
		Trees_din <= x"00361041";
		wait for Clk_period;
		Addr <=  "00001111100111";
		Trees_din <= x"0018d034";
		wait for Clk_period;
		Addr <=  "00001111101000";
		Trees_din <= x"0113e920";
		wait for Clk_period;
		Addr <=  "00001111101001";
		Trees_din <= x"0c03cc10";
		wait for Clk_period;
		Addr <=  "00001111101010";
		Trees_din <= x"07005608";
		wait for Clk_period;
		Addr <=  "00001111101011";
		Trees_din <= x"09005104";
		wait for Clk_period;
		Addr <=  "00001111101100";
		Trees_din <= x"00291041";
		wait for Clk_period;
		Addr <=  "00001111101101";
		Trees_din <= x"ffe71041";
		wait for Clk_period;
		Addr <=  "00001111101110";
		Trees_din <= x"07005704";
		wait for Clk_period;
		Addr <=  "00001111101111";
		Trees_din <= x"00681041";
		wait for Clk_period;
		Addr <=  "00001111110000";
		Trees_din <= x"00131041";
		wait for Clk_period;
		Addr <=  "00001111110001";
		Trees_din <= x"19008d08";
		wait for Clk_period;
		Addr <=  "00001111110010";
		Trees_din <= x"0afb2604";
		wait for Clk_period;
		Addr <=  "00001111110011";
		Trees_din <= x"00171041";
		wait for Clk_period;
		Addr <=  "00001111110100";
		Trees_din <= x"00e61041";
		wait for Clk_period;
		Addr <=  "00001111110101";
		Trees_din <= x"08019304";
		wait for Clk_period;
		Addr <=  "00001111110110";
		Trees_din <= x"ff9a1041";
		wait for Clk_period;
		Addr <=  "00001111110111";
		Trees_din <= x"00711041";
		wait for Clk_period;
		Addr <=  "00001111111000";
		Trees_din <= x"000f0708";
		wait for Clk_period;
		Addr <=  "00001111111001";
		Trees_din <= x"0209bd04";
		wait for Clk_period;
		Addr <=  "00001111111010";
		Trees_din <= x"009c1041";
		wait for Clk_period;
		Addr <=  "00001111111011";
		Trees_din <= x"00141041";
		wait for Clk_period;
		Addr <=  "00001111111100";
		Trees_din <= x"0ef98004";
		wait for Clk_period;
		Addr <=  "00001111111101";
		Trees_din <= x"ff7e1041";
		wait for Clk_period;
		Addr <=  "00001111111110";
		Trees_din <= x"1d005104";
		wait for Clk_period;
		Addr <=  "00001111111111";
		Trees_din <= x"00661041";
		wait for Clk_period;
		Addr <=  "00010000000000";
		Trees_din <= x"ffcf1041";
		wait for Clk_period;
		Addr <=  "00010000000001";
		Trees_din <= x"010ed010";
		wait for Clk_period;
		Addr <=  "00010000000010";
		Trees_din <= x"0f03d408";
		wait for Clk_period;
		Addr <=  "00010000000011";
		Trees_din <= x"0e043e04";
		wait for Clk_period;
		Addr <=  "00010000000100";
		Trees_din <= x"ff6b1041";
		wait for Clk_period;
		Addr <=  "00010000000101";
		Trees_din <= x"00321041";
		wait for Clk_period;
		Addr <=  "00010000000110";
		Trees_din <= x"18003f04";
		wait for Clk_period;
		Addr <=  "00010000000111";
		Trees_din <= x"00df1041";
		wait for Clk_period;
		Addr <=  "00010000001000";
		Trees_din <= x"ff931041";
		wait for Clk_period;
		Addr <=  "00010000001001";
		Trees_din <= x"1900980c";
		wait for Clk_period;
		Addr <=  "00010000001010";
		Trees_din <= x"1a00b704";
		wait for Clk_period;
		Addr <=  "00010000001011";
		Trees_din <= x"ffa41041";
		wait for Clk_period;
		Addr <=  "00010000001100";
		Trees_din <= x"0201e304";
		wait for Clk_period;
		Addr <=  "00010000001101";
		Trees_din <= x"00e01041";
		wait for Clk_period;
		Addr <=  "00010000001110";
		Trees_din <= x"00271041";
		wait for Clk_period;
		Addr <=  "00010000001111";
		Trees_din <= x"ff8e1041";
		wait for Clk_period;
		Addr <=  "00010000010000";
		Trees_din <= x"01017520";
		wait for Clk_period;
		Addr <=  "00010000010001";
		Trees_din <= x"0f03e610";
		wait for Clk_period;
		Addr <=  "00010000010010";
		Trees_din <= x"07005e0c";
		wait for Clk_period;
		Addr <=  "00010000010011";
		Trees_din <= x"0af83808";
		wait for Clk_period;
		Addr <=  "00010000010100";
		Trees_din <= x"0800e204";
		wait for Clk_period;
		Addr <=  "00010000010101";
		Trees_din <= x"ff7f10f5";
		wait for Clk_period;
		Addr <=  "00010000010110";
		Trees_din <= x"003e10f5";
		wait for Clk_period;
		Addr <=  "00010000010111";
		Trees_din <= x"ff6810f5";
		wait for Clk_period;
		Addr <=  "00010000011000";
		Trees_din <= x"000c10f5";
		wait for Clk_period;
		Addr <=  "00010000011001";
		Trees_din <= x"1101220c";
		wait for Clk_period;
		Addr <=  "00010000011010";
		Trees_din <= x"02009004";
		wait for Clk_period;
		Addr <=  "00010000011011";
		Trees_din <= x"ffb110f5";
		wait for Clk_period;
		Addr <=  "00010000011100";
		Trees_din <= x"0302da04";
		wait for Clk_period;
		Addr <=  "00010000011101";
		Trees_din <= x"001210f5";
		wait for Clk_period;
		Addr <=  "00010000011110";
		Trees_din <= x"00af10f5";
		wait for Clk_period;
		Addr <=  "00010000011111";
		Trees_din <= x"ff8d10f5";
		wait for Clk_period;
		Addr <=  "00010000100000";
		Trees_din <= x"001fa434";
		wait for Clk_period;
		Addr <=  "00010000100001";
		Trees_din <= x"01159320";
		wait for Clk_period;
		Addr <=  "00010000100010";
		Trees_din <= x"010a4210";
		wait for Clk_period;
		Addr <=  "00010000100011";
		Trees_din <= x"0b04a108";
		wait for Clk_period;
		Addr <=  "00010000100100";
		Trees_din <= x"18004c04";
		wait for Clk_period;
		Addr <=  "00010000100101";
		Trees_din <= x"001c10f5";
		wait for Clk_period;
		Addr <=  "00010000100110";
		Trees_din <= x"ffbd10f5";
		wait for Clk_period;
		Addr <=  "00010000100111";
		Trees_din <= x"15009804";
		wait for Clk_period;
		Addr <=  "00010000101000";
		Trees_din <= x"000410f5";
		wait for Clk_period;
		Addr <=  "00010000101001";
		Trees_din <= x"ff8610f5";
		wait for Clk_period;
		Addr <=  "00010000101010";
		Trees_din <= x"05fa4108";
		wait for Clk_period;
		Addr <=  "00010000101011";
		Trees_din <= x"0c02dd04";
		wait for Clk_period;
		Addr <=  "00010000101100";
		Trees_din <= x"fff510f5";
		wait for Clk_period;
		Addr <=  "00010000101101";
		Trees_din <= x"004510f5";
		wait for Clk_period;
		Addr <=  "00010000101110";
		Trees_din <= x"11046d04";
		wait for Clk_period;
		Addr <=  "00010000101111";
		Trees_din <= x"004b10f5";
		wait for Clk_period;
		Addr <=  "00010000110000";
		Trees_din <= x"ffc210f5";
		wait for Clk_period;
		Addr <=  "00010000110001";
		Trees_din <= x"0b046008";
		wait for Clk_period;
		Addr <=  "00010000110010";
		Trees_din <= x"1203bc04";
		wait for Clk_period;
		Addr <=  "00010000110011";
		Trees_din <= x"009810f5";
		wait for Clk_period;
		Addr <=  "00010000110100";
		Trees_din <= x"002e10f5";
		wait for Clk_period;
		Addr <=  "00010000110101";
		Trees_din <= x"00132408";
		wait for Clk_period;
		Addr <=  "00010000110110";
		Trees_din <= x"1c002804";
		wait for Clk_period;
		Addr <=  "00010000110111";
		Trees_din <= x"000d10f5";
		wait for Clk_period;
		Addr <=  "00010000111000";
		Trees_din <= x"007910f5";
		wait for Clk_period;
		Addr <=  "00010000111001";
		Trees_din <= x"ffab10f5";
		wait for Clk_period;
		Addr <=  "00010000111010";
		Trees_din <= x"1f000104";
		wait for Clk_period;
		Addr <=  "00010000111011";
		Trees_din <= x"ff7010f5";
		wait for Clk_period;
		Addr <=  "00010000111100";
		Trees_din <= x"004b10f5";
		wait for Clk_period;
		Addr <=  "00010000111101";
		Trees_din <= x"0101751c";
		wait for Clk_period;
		Addr <=  "00010000111110";
		Trees_din <= x"0f03e610";
		wait for Clk_period;
		Addr <=  "00010000111111";
		Trees_din <= x"07005e0c";
		wait for Clk_period;
		Addr <=  "00010001000000";
		Trees_din <= x"0af83808";
		wait for Clk_period;
		Addr <=  "00010001000001";
		Trees_din <= x"0800e204";
		wait for Clk_period;
		Addr <=  "00010001000010";
		Trees_din <= x"ff8411a1";
		wait for Clk_period;
		Addr <=  "00010001000011";
		Trees_din <= x"004111a1";
		wait for Clk_period;
		Addr <=  "00010001000100";
		Trees_din <= x"ff6a11a1";
		wait for Clk_period;
		Addr <=  "00010001000101";
		Trees_din <= x"001311a1";
		wait for Clk_period;
		Addr <=  "00010001000110";
		Trees_din <= x"11012208";
		wait for Clk_period;
		Addr <=  "00010001000111";
		Trees_din <= x"07005a04";
		wait for Clk_period;
		Addr <=  "00010001001000";
		Trees_din <= x"ffed11a1";
		wait for Clk_period;
		Addr <=  "00010001001001";
		Trees_din <= x"007f11a1";
		wait for Clk_period;
		Addr <=  "00010001001010";
		Trees_din <= x"ff9411a1";
		wait for Clk_period;
		Addr <=  "00010001001011";
		Trees_din <= x"001fa434";
		wait for Clk_period;
		Addr <=  "00010001001100";
		Trees_din <= x"01159320";
		wait for Clk_period;
		Addr <=  "00010001001101";
		Trees_din <= x"05fcb210";
		wait for Clk_period;
		Addr <=  "00010001001110";
		Trees_din <= x"05fc9d08";
		wait for Clk_period;
		Addr <=  "00010001001111";
		Trees_din <= x"1900a404";
		wait for Clk_period;
		Addr <=  "00010001010000";
		Trees_din <= x"002011a1";
		wait for Clk_period;
		Addr <=  "00010001010001";
		Trees_din <= x"fff111a1";
		wait for Clk_period;
		Addr <=  "00010001010010";
		Trees_din <= x"09005204";
		wait for Clk_period;
		Addr <=  "00010001010011";
		Trees_din <= x"ff9311a1";
		wait for Clk_period;
		Addr <=  "00010001010100";
		Trees_din <= x"011411a1";
		wait for Clk_period;
		Addr <=  "00010001010101";
		Trees_din <= x"1b003a08";
		wait for Clk_period;
		Addr <=  "00010001010110";
		Trees_din <= x"0201e304";
		wait for Clk_period;
		Addr <=  "00010001010111";
		Trees_din <= x"005f11a1";
		wait for Clk_period;
		Addr <=  "00010001011000";
		Trees_din <= x"ffd611a1";
		wait for Clk_period;
		Addr <=  "00010001011001";
		Trees_din <= x"05fe1904";
		wait for Clk_period;
		Addr <=  "00010001011010";
		Trees_din <= x"ff7e11a1";
		wait for Clk_period;
		Addr <=  "00010001011011";
		Trees_din <= x"000811a1";
		wait for Clk_period;
		Addr <=  "00010001011100";
		Trees_din <= x"0b046008";
		wait for Clk_period;
		Addr <=  "00010001011101";
		Trees_din <= x"10fa6104";
		wait for Clk_period;
		Addr <=  "00010001011110";
		Trees_din <= x"002d11a1";
		wait for Clk_period;
		Addr <=  "00010001011111";
		Trees_din <= x"009411a1";
		wait for Clk_period;
		Addr <=  "00010001100000";
		Trees_din <= x"15008904";
		wait for Clk_period;
		Addr <=  "00010001100001";
		Trees_din <= x"ffb411a1";
		wait for Clk_period;
		Addr <=  "00010001100010";
		Trees_din <= x"1500a804";
		wait for Clk_period;
		Addr <=  "00010001100011";
		Trees_din <= x"007411a1";
		wait for Clk_period;
		Addr <=  "00010001100100";
		Trees_din <= x"000a11a1";
		wait for Clk_period;
		Addr <=  "00010001100101";
		Trees_din <= x"1900ab04";
		wait for Clk_period;
		Addr <=  "00010001100110";
		Trees_din <= x"ff7311a1";
		wait for Clk_period;
		Addr <=  "00010001100111";
		Trees_din <= x"002b11a1";
		wait for Clk_period;
		Addr <=  "00010001101000";
		Trees_din <= x"01017518";
		wait for Clk_period;
		Addr <=  "00010001101001";
		Trees_din <= x"15008b0c";
		wait for Clk_period;
		Addr <=  "00010001101010";
		Trees_din <= x"15008908";
		wait for Clk_period;
		Addr <=  "00010001101011";
		Trees_din <= x"1403f904";
		wait for Clk_period;
		Addr <=  "00010001101100";
		Trees_din <= x"ff79123d";
		wait for Clk_period;
		Addr <=  "00010001101101";
		Trees_din <= x"0047123d";
		wait for Clk_period;
		Addr <=  "00010001101110";
		Trees_din <= x"00ba123d";
		wait for Clk_period;
		Addr <=  "00010001101111";
		Trees_din <= x"10f7fb08";
		wait for Clk_period;
		Addr <=  "00010001110000";
		Trees_din <= x"17001204";
		wait for Clk_period;
		Addr <=  "00010001110001";
		Trees_din <= x"0028123d";
		wait for Clk_period;
		Addr <=  "00010001110010";
		Trees_din <= x"ffa3123d";
		wait for Clk_period;
		Addr <=  "00010001110011";
		Trees_din <= x"ff6b123d";
		wait for Clk_period;
		Addr <=  "00010001110100";
		Trees_din <= x"00229234";
		wait for Clk_period;
		Addr <=  "00010001110101";
		Trees_din <= x"01159320";
		wait for Clk_period;
		Addr <=  "00010001110110";
		Trees_din <= x"0f00c310";
		wait for Clk_period;
		Addr <=  "00010001110111";
		Trees_din <= x"01096908";
		wait for Clk_period;
		Addr <=  "00010001111000";
		Trees_din <= x"07005d04";
		wait for Clk_period;
		Addr <=  "00010001111001";
		Trees_din <= x"ffca123d";
		wait for Clk_period;
		Addr <=  "00010001111010";
		Trees_din <= x"00a0123d";
		wait for Clk_period;
		Addr <=  "00010001111011";
		Trees_din <= x"1400ef04";
		wait for Clk_period;
		Addr <=  "00010001111100";
		Trees_din <= x"002c123d";
		wait for Clk_period;
		Addr <=  "00010001111101";
		Trees_din <= x"ffda123d";
		wait for Clk_period;
		Addr <=  "00010001111110";
		Trees_din <= x"14027c08";
		wait for Clk_period;
		Addr <=  "00010001111111";
		Trees_din <= x"03fbf604";
		wait for Clk_period;
		Addr <=  "00010010000000";
		Trees_din <= x"001c123d";
		wait for Clk_period;
		Addr <=  "00010010000001";
		Trees_din <= x"006e123d";
		wait for Clk_period;
		Addr <=  "00010010000010";
		Trees_din <= x"12028704";
		wait for Clk_period;
		Addr <=  "00010010000011";
		Trees_din <= x"0019123d";
		wait for Clk_period;
		Addr <=  "00010010000100";
		Trees_din <= x"ffbc123d";
		wait for Clk_period;
		Addr <=  "00010010000101";
		Trees_din <= x"0b046008";
		wait for Clk_period;
		Addr <=  "00010010000110";
		Trees_din <= x"1c002604";
		wait for Clk_period;
		Addr <=  "00010010000111";
		Trees_din <= x"0017123d";
		wait for Clk_period;
		Addr <=  "00010010001000";
		Trees_din <= x"008c123d";
		wait for Clk_period;
		Addr <=  "00010010001001";
		Trees_din <= x"00132408";
		wait for Clk_period;
		Addr <=  "00010010001010";
		Trees_din <= x"0afa1a04";
		wait for Clk_period;
		Addr <=  "00010010001011";
		Trees_din <= x"000a123d";
		wait for Clk_period;
		Addr <=  "00010010001100";
		Trees_din <= x"006d123d";
		wait for Clk_period;
		Addr <=  "00010010001101";
		Trees_din <= x"ffba123d";
		wait for Clk_period;
		Addr <=  "00010010001110";
		Trees_din <= x"ff7b123d";
		wait for Clk_period;
		Addr <=  "00010010001111";
		Trees_din <= x"01017518";
		wait for Clk_period;
		Addr <=  "00010010010000";
		Trees_din <= x"15008b0c";
		wait for Clk_period;
		Addr <=  "00010010010001";
		Trees_din <= x"15008908";
		wait for Clk_period;
		Addr <=  "00010010010010";
		Trees_din <= x"1403f904";
		wait for Clk_period;
		Addr <=  "00010010010011";
		Trees_din <= x"ff7d1309";
		wait for Clk_period;
		Addr <=  "00010010010100";
		Trees_din <= x"00401309";
		wait for Clk_period;
		Addr <=  "00010010010101";
		Trees_din <= x"00a01309";
		wait for Clk_period;
		Addr <=  "00010010010110";
		Trees_din <= x"06f35808";
		wait for Clk_period;
		Addr <=  "00010010010111";
		Trees_din <= x"02027c04";
		wait for Clk_period;
		Addr <=  "00010010011000";
		Trees_din <= x"00251309";
		wait for Clk_period;
		Addr <=  "00010010011001";
		Trees_din <= x"ffac1309";
		wait for Clk_period;
		Addr <=  "00010010011010";
		Trees_din <= x"ff6d1309";
		wait for Clk_period;
		Addr <=  "00010010011011";
		Trees_din <= x"0115933c";
		wait for Clk_period;
		Addr <=  "00010010011100";
		Trees_din <= x"04f69f1c";
		wait for Clk_period;
		Addr <=  "00010010011101";
		Trees_din <= x"03fc5310";
		wait for Clk_period;
		Addr <=  "00010010011110";
		Trees_din <= x"1f000208";
		wait for Clk_period;
		Addr <=  "00010010011111";
		Trees_din <= x"010bb604";
		wait for Clk_period;
		Addr <=  "00010010100000";
		Trees_din <= x"ff711309";
		wait for Clk_period;
		Addr <=  "00010010100001";
		Trees_din <= x"ffe71309";
		wait for Clk_period;
		Addr <=  "00010010100010";
		Trees_din <= x"08007b04";
		wait for Clk_period;
		Addr <=  "00010010100011";
		Trees_din <= x"01121309";
		wait for Clk_period;
		Addr <=  "00010010100100";
		Trees_din <= x"ffe01309";
		wait for Clk_period;
		Addr <=  "00010010100101";
		Trees_din <= x"05f94a08";
		wait for Clk_period;
		Addr <=  "00010010100110";
		Trees_din <= x"01092404";
		wait for Clk_period;
		Addr <=  "00010010100111";
		Trees_din <= x"ff911309";
		wait for Clk_period;
		Addr <=  "00010010101000";
		Trees_din <= x"00601309";
		wait for Clk_period;
		Addr <=  "00010010101001";
		Trees_din <= x"01291309";
		wait for Clk_period;
		Addr <=  "00010010101010";
		Trees_din <= x"0c001910";
		wait for Clk_period;
		Addr <=  "00010010101011";
		Trees_din <= x"0e008808";
		wait for Clk_period;
		Addr <=  "00010010101100";
		Trees_din <= x"0b040404";
		wait for Clk_period;
		Addr <=  "00010010101101";
		Trees_din <= x"01391309";
		wait for Clk_period;
		Addr <=  "00010010101110";
		Trees_din <= x"00391309";
		wait for Clk_period;
		Addr <=  "00010010101111";
		Trees_din <= x"03fb7404";
		wait for Clk_period;
		Addr <=  "00010010110000";
		Trees_din <= x"fffb1309";
		wait for Clk_period;
		Addr <=  "00010010110001";
		Trees_din <= x"ff8b1309";
		wait for Clk_period;
		Addr <=  "00010010110010";
		Trees_din <= x"1603f908";
		wait for Clk_period;
		Addr <=  "00010010110011";
		Trees_din <= x"04f6f504";
		wait for Clk_period;
		Addr <=  "00010010110100";
		Trees_din <= x"009d1309";
		wait for Clk_period;
		Addr <=  "00010010110101";
		Trees_din <= x"00121309";
		wait for Clk_period;
		Addr <=  "00010010110110";
		Trees_din <= x"0a03a304";
		wait for Clk_period;
		Addr <=  "00010010110111";
		Trees_din <= x"ffb41309";
		wait for Clk_period;
		Addr <=  "00010010111000";
		Trees_din <= x"007d1309";
		wait for Clk_period;
		Addr <=  "00010010111001";
		Trees_din <= x"0013bd08";
		wait for Clk_period;
		Addr <=  "00010010111010";
		Trees_din <= x"02080c04";
		wait for Clk_period;
		Addr <=  "00010010111011";
		Trees_din <= x"008f1309";
		wait for Clk_period;
		Addr <=  "00010010111100";
		Trees_din <= x"001a1309";
		wait for Clk_period;
		Addr <=  "00010010111101";
		Trees_din <= x"15008904";
		wait for Clk_period;
		Addr <=  "00010010111110";
		Trees_din <= x"ffbf1309";
		wait for Clk_period;
		Addr <=  "00010010111111";
		Trees_din <= x"0d010904";
		wait for Clk_period;
		Addr <=  "00010011000000";
		Trees_din <= x"fff71309";
		wait for Clk_period;
		Addr <=  "00010011000001";
		Trees_din <= x"007f1309";
		wait for Clk_period;
		Addr <=  "00010011000010";
		Trees_din <= x"01017518";
		wait for Clk_period;
		Addr <=  "00010011000011";
		Trees_din <= x"15008b10";
		wait for Clk_period;
		Addr <=  "00010011000100";
		Trees_din <= x"15008908";
		wait for Clk_period;
		Addr <=  "00010011000101";
		Trees_din <= x"1403f904";
		wait for Clk_period;
		Addr <=  "00010011000110";
		Trees_din <= x"ff8113cd";
		wait for Clk_period;
		Addr <=  "00010011000111";
		Trees_din <= x"003a13cd";
		wait for Clk_period;
		Addr <=  "00010011001000";
		Trees_din <= x"0d027504";
		wait for Clk_period;
		Addr <=  "00010011001001";
		Trees_din <= x"ffff13cd";
		wait for Clk_period;
		Addr <=  "00010011001010";
		Trees_din <= x"00d013cd";
		wait for Clk_period;
		Addr <=  "00010011001011";
		Trees_din <= x"10f7fb04";
		wait for Clk_period;
		Addr <=  "00010011001100";
		Trees_din <= x"ffe713cd";
		wait for Clk_period;
		Addr <=  "00010011001101";
		Trees_din <= x"ff6e13cd";
		wait for Clk_period;
		Addr <=  "00010011001110";
		Trees_din <= x"01159338";
		wait for Clk_period;
		Addr <=  "00010011001111";
		Trees_din <= x"13fa0b18";
		wait for Clk_period;
		Addr <=  "00010011010000";
		Trees_din <= x"0a012808";
		wait for Clk_period;
		Addr <=  "00010011010001";
		Trees_din <= x"14007d04";
		wait for Clk_period;
		Addr <=  "00010011010010";
		Trees_din <= x"001313cd";
		wait for Clk_period;
		Addr <=  "00010011010011";
		Trees_din <= x"ff5513cd";
		wait for Clk_period;
		Addr <=  "00010011010100";
		Trees_din <= x"05f8c108";
		wait for Clk_period;
		Addr <=  "00010011010101";
		Trees_din <= x"19007d04";
		wait for Clk_period;
		Addr <=  "00010011010110";
		Trees_din <= x"007e13cd";
		wait for Clk_period;
		Addr <=  "00010011010111";
		Trees_din <= x"ff8913cd";
		wait for Clk_period;
		Addr <=  "00010011011000";
		Trees_din <= x"0efdf804";
		wait for Clk_period;
		Addr <=  "00010011011001";
		Trees_din <= x"003413cd";
		wait for Clk_period;
		Addr <=  "00010011011010";
		Trees_din <= x"ffd013cd";
		wait for Clk_period;
		Addr <=  "00010011011011";
		Trees_din <= x"1f000010";
		wait for Clk_period;
		Addr <=  "00010011011100";
		Trees_din <= x"04f5dd08";
		wait for Clk_period;
		Addr <=  "00010011011101";
		Trees_din <= x"0f000a04";
		wait for Clk_period;
		Addr <=  "00010011011110";
		Trees_din <= x"005e13cd";
		wait for Clk_period;
		Addr <=  "00010011011111";
		Trees_din <= x"ffa713cd";
		wait for Clk_period;
		Addr <=  "00010011100000";
		Trees_din <= x"0802a504";
		wait for Clk_period;
		Addr <=  "00010011100001";
		Trees_din <= x"001813cd";
		wait for Clk_period;
		Addr <=  "00010011100010";
		Trees_din <= x"006513cd";
		wait for Clk_period;
		Addr <=  "00010011100011";
		Trees_din <= x"0b04ee08";
		wait for Clk_period;
		Addr <=  "00010011100100";
		Trees_din <= x"1a00ba04";
		wait for Clk_period;
		Addr <=  "00010011100101";
		Trees_din <= x"007f13cd";
		wait for Clk_period;
		Addr <=  "00010011100110";
		Trees_din <= x"ff9b13cd";
		wait for Clk_period;
		Addr <=  "00010011100111";
		Trees_din <= x"0c02b104";
		wait for Clk_period;
		Addr <=  "00010011101000";
		Trees_din <= x"00e313cd";
		wait for Clk_period;
		Addr <=  "00010011101001";
		Trees_din <= x"ffc313cd";
		wait for Clk_period;
		Addr <=  "00010011101010";
		Trees_din <= x"0013bd08";
		wait for Clk_period;
		Addr <=  "00010011101011";
		Trees_din <= x"02080c04";
		wait for Clk_period;
		Addr <=  "00010011101100";
		Trees_din <= x"008b13cd";
		wait for Clk_period;
		Addr <=  "00010011101101";
		Trees_din <= x"001613cd";
		wait for Clk_period;
		Addr <=  "00010011101110";
		Trees_din <= x"15008904";
		wait for Clk_period;
		Addr <=  "00010011101111";
		Trees_din <= x"ffc613cd";
		wait for Clk_period;
		Addr <=  "00010011110000";
		Trees_din <= x"0d010904";
		wait for Clk_period;
		Addr <=  "00010011110001";
		Trees_din <= x"fffa13cd";
		wait for Clk_period;
		Addr <=  "00010011110010";
		Trees_din <= x"007713cd";
		wait for Clk_period;
		Addr <=  "00010011110011";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00010011110100";
		Trees_din <= x"01017518";
		wait for Clk_period;
		Addr <=  "00010011110101";
		Trees_din <= x"15008b10";
		wait for Clk_period;
		Addr <=  "00010011110110";
		Trees_din <= x"18004908";
		wait for Clk_period;
		Addr <=  "00010011110111";
		Trees_din <= x"02025f04";
		wait for Clk_period;
		Addr <=  "00010011111000";
		Trees_din <= x"fff114b5";
		wait for Clk_period;
		Addr <=  "00010011111001";
		Trees_din <= x"00dc14b5";
		wait for Clk_period;
		Addr <=  "00010011111010";
		Trees_din <= x"09005c04";
		wait for Clk_period;
		Addr <=  "00010011111011";
		Trees_din <= x"ff8414b5";
		wait for Clk_period;
		Addr <=  "00010011111100";
		Trees_din <= x"003314b5";
		wait for Clk_period;
		Addr <=  "00010011111101";
		Trees_din <= x"0f03e604";
		wait for Clk_period;
		Addr <=  "00010011111110";
		Trees_din <= x"ff7014b5";
		wait for Clk_period;
		Addr <=  "00010011111111";
		Trees_din <= x"fff014b5";
		wait for Clk_period;
		Addr <=  "00010100000000";
		Trees_din <= x"0113e934";
		wait for Clk_period;
		Addr <=  "00010100000001";
		Trees_din <= x"0c003218";
		wait for Clk_period;
		Addr <=  "00010100000010";
		Trees_din <= x"05fb4a0c";
		wait for Clk_period;
		Addr <=  "00010100000011";
		Trees_din <= x"0d00c408";
		wait for Clk_period;
		Addr <=  "00010100000100";
		Trees_din <= x"18004c04";
		wait for Clk_period;
		Addr <=  "00010100000101";
		Trees_din <= x"00dc14b5";
		wait for Clk_period;
		Addr <=  "00010100000110";
		Trees_din <= x"000214b5";
		wait for Clk_period;
		Addr <=  "00010100000111";
		Trees_din <= x"ffaf14b5";
		wait for Clk_period;
		Addr <=  "00010100001000";
		Trees_din <= x"04fd9804";
		wait for Clk_period;
		Addr <=  "00010100001001";
		Trees_din <= x"ff6c14b5";
		wait for Clk_period;
		Addr <=  "00010100001010";
		Trees_din <= x"03fbbc04";
		wait for Clk_period;
		Addr <=  "00010100001011";
		Trees_din <= x"00be14b5";
		wait for Clk_period;
		Addr <=  "00010100001100";
		Trees_din <= x"ffc614b5";
		wait for Clk_period;
		Addr <=  "00010100001101";
		Trees_din <= x"1603fa10";
		wait for Clk_period;
		Addr <=  "00010100001110";
		Trees_din <= x"0d000508";
		wait for Clk_period;
		Addr <=  "00010100001111";
		Trees_din <= x"1d004804";
		wait for Clk_period;
		Addr <=  "00010100010000";
		Trees_din <= x"ff8114b5";
		wait for Clk_period;
		Addr <=  "00010100010001";
		Trees_din <= x"000d14b5";
		wait for Clk_period;
		Addr <=  "00010100010010";
		Trees_din <= x"07005604";
		wait for Clk_period;
		Addr <=  "00010100010011";
		Trees_din <= x"fffc14b5";
		wait for Clk_period;
		Addr <=  "00010100010100";
		Trees_din <= x"001e14b5";
		wait for Clk_period;
		Addr <=  "00010100010101";
		Trees_din <= x"19009b08";
		wait for Clk_period;
		Addr <=  "00010100010110";
		Trees_din <= x"1a00bd04";
		wait for Clk_period;
		Addr <=  "00010100010111";
		Trees_din <= x"ff6f14b5";
		wait for Clk_period;
		Addr <=  "00010100011000";
		Trees_din <= x"005114b5";
		wait for Clk_period;
		Addr <=  "00010100011001";
		Trees_din <= x"ff5314b5";
		wait for Clk_period;
		Addr <=  "00010100011010";
		Trees_din <= x"1a00e018";
		wait for Clk_period;
		Addr <=  "00010100011011";
		Trees_din <= x"00148708";
		wait for Clk_period;
		Addr <=  "00010100011100";
		Trees_din <= x"1d005604";
		wait for Clk_period;
		Addr <=  "00010100011101";
		Trees_din <= x"009514b5";
		wait for Clk_period;
		Addr <=  "00010100011110";
		Trees_din <= x"000714b5";
		wait for Clk_period;
		Addr <=  "00010100011111";
		Trees_din <= x"16018508";
		wait for Clk_period;
		Addr <=  "00010100100000";
		Trees_din <= x"11028a04";
		wait for Clk_period;
		Addr <=  "00010100100001";
		Trees_din <= x"ff9d14b5";
		wait for Clk_period;
		Addr <=  "00010100100010";
		Trees_din <= x"002314b5";
		wait for Clk_period;
		Addr <=  "00010100100011";
		Trees_din <= x"1c003704";
		wait for Clk_period;
		Addr <=  "00010100100100";
		Trees_din <= x"001014b5";
		wait for Clk_period;
		Addr <=  "00010100100101";
		Trees_din <= x"006814b5";
		wait for Clk_period;
		Addr <=  "00010100100110";
		Trees_din <= x"01159308";
		wait for Clk_period;
		Addr <=  "00010100100111";
		Trees_din <= x"0f00a604";
		wait for Clk_period;
		Addr <=  "00010100101000";
		Trees_din <= x"fff614b5";
		wait for Clk_period;
		Addr <=  "00010100101001";
		Trees_din <= x"ff6f14b5";
		wait for Clk_period;
		Addr <=  "00010100101010";
		Trees_din <= x"0afd0204";
		wait for Clk_period;
		Addr <=  "00010100101011";
		Trees_din <= x"ffe514b5";
		wait for Clk_period;
		Addr <=  "00010100101100";
		Trees_din <= x"006d14b5";
		wait for Clk_period;
		Addr <=  "00010100101101";
		Trees_din <= x"01fe6a04";
		wait for Clk_period;
		Addr <=  "00010100101110";
		Trees_din <= x"ff761589";
		wait for Clk_period;
		Addr <=  "00010100101111";
		Trees_din <= x"010a4234";
		wait for Clk_period;
		Addr <=  "00010100110000";
		Trees_din <= x"0b04a118";
		wait for Clk_period;
		Addr <=  "00010100110001";
		Trees_din <= x"04f56808";
		wait for Clk_period;
		Addr <=  "00010100110010";
		Trees_din <= x"10055d04";
		wait for Clk_period;
		Addr <=  "00010100110011";
		Trees_din <= x"ff6d1589";
		wait for Clk_period;
		Addr <=  "00010100110100";
		Trees_din <= x"00261589";
		wait for Clk_period;
		Addr <=  "00010100110101";
		Trees_din <= x"12038808";
		wait for Clk_period;
		Addr <=  "00010100110110";
		Trees_din <= x"1f000004";
		wait for Clk_period;
		Addr <=  "00010100110111";
		Trees_din <= x"00241589";
		wait for Clk_period;
		Addr <=  "00010100111000";
		Trees_din <= x"ffb21589";
		wait for Clk_period;
		Addr <=  "00010100111001";
		Trees_din <= x"0802c204";
		wait for Clk_period;
		Addr <=  "00010100111010";
		Trees_din <= x"ff951589";
		wait for Clk_period;
		Addr <=  "00010100111011";
		Trees_din <= x"00911589";
		wait for Clk_period;
		Addr <=  "00010100111100";
		Trees_din <= x"0e003410";
		wait for Clk_period;
		Addr <=  "00010100111101";
		Trees_din <= x"13ff1308";
		wait for Clk_period;
		Addr <=  "00010100111110";
		Trees_din <= x"1100a204";
		wait for Clk_period;
		Addr <=  "00010100111111";
		Trees_din <= x"ffc21589";
		wait for Clk_period;
		Addr <=  "00010101000000";
		Trees_din <= x"00a91589";
		wait for Clk_period;
		Addr <=  "00010101000001";
		Trees_din <= x"11fda704";
		wait for Clk_period;
		Addr <=  "00010101000010";
		Trees_din <= x"fff41589";
		wait for Clk_period;
		Addr <=  "00010101000011";
		Trees_din <= x"01371589";
		wait for Clk_period;
		Addr <=  "00010101000100";
		Trees_din <= x"06fb2908";
		wait for Clk_period;
		Addr <=  "00010101000101";
		Trees_din <= x"07004d04";
		wait for Clk_period;
		Addr <=  "00010101000110";
		Trees_din <= x"00211589";
		wait for Clk_period;
		Addr <=  "00010101000111";
		Trees_din <= x"ff511589";
		wait for Clk_period;
		Addr <=  "00010101001000";
		Trees_din <= x"003a1589";
		wait for Clk_period;
		Addr <=  "00010101001001";
		Trees_din <= x"05fb0f20";
		wait for Clk_period;
		Addr <=  "00010101001010";
		Trees_din <= x"09005810";
		wait for Clk_period;
		Addr <=  "00010101001011";
		Trees_din <= x"06f68b08";
		wait for Clk_period;
		Addr <=  "00010101001100";
		Trees_din <= x"0c011c04";
		wait for Clk_period;
		Addr <=  "00010101001101";
		Trees_din <= x"ffcc1589";
		wait for Clk_period;
		Addr <=  "00010101001110";
		Trees_din <= x"001d1589";
		wait for Clk_period;
		Addr <=  "00010101001111";
		Trees_din <= x"11028704";
		wait for Clk_period;
		Addr <=  "00010101010000";
		Trees_din <= x"006b1589";
		wait for Clk_period;
		Addr <=  "00010101010001";
		Trees_din <= x"ffe71589";
		wait for Clk_period;
		Addr <=  "00010101010010";
		Trees_din <= x"07005b08";
		wait for Clk_period;
		Addr <=  "00010101010011";
		Trees_din <= x"02ff8604";
		wait for Clk_period;
		Addr <=  "00010101010100";
		Trees_din <= x"00841589";
		wait for Clk_period;
		Addr <=  "00010101010101";
		Trees_din <= x"ffa01589";
		wait for Clk_period;
		Addr <=  "00010101010110";
		Trees_din <= x"1d004f04";
		wait for Clk_period;
		Addr <=  "00010101010111";
		Trees_din <= x"00901589";
		wait for Clk_period;
		Addr <=  "00010101011000";
		Trees_din <= x"ffb41589";
		wait for Clk_period;
		Addr <=  "00010101011001";
		Trees_din <= x"14001304";
		wait for Clk_period;
		Addr <=  "00010101011010";
		Trees_din <= x"ff581589";
		wait for Clk_period;
		Addr <=  "00010101011011";
		Trees_din <= x"07005508";
		wait for Clk_period;
		Addr <=  "00010101011100";
		Trees_din <= x"19008a04";
		wait for Clk_period;
		Addr <=  "00010101011101";
		Trees_din <= x"00b01589";
		wait for Clk_period;
		Addr <=  "00010101011110";
		Trees_din <= x"ffc91589";
		wait for Clk_period;
		Addr <=  "00010101011111";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00010101100000";
		Trees_din <= x"00a01589";
		wait for Clk_period;
		Addr <=  "00010101100001";
		Trees_din <= x"000c1589";
		wait for Clk_period;
		Addr <=  "00010101100010";
		Trees_din <= x"01fe6a04";
		wait for Clk_period;
		Addr <=  "00010101100011";
		Trees_din <= x"ff781615";
		wait for Clk_period;
		Addr <=  "00010101100100";
		Trees_din <= x"01159334";
		wait for Clk_period;
		Addr <=  "00010101100101";
		Trees_din <= x"2004001c";
		wait for Clk_period;
		Addr <=  "00010101100110";
		Trees_din <= x"05f9a40c";
		wait for Clk_period;
		Addr <=  "00010101100111";
		Trees_din <= x"19009e08";
		wait for Clk_period;
		Addr <=  "00010101101000";
		Trees_din <= x"04f72f04";
		wait for Clk_period;
		Addr <=  "00010101101001";
		Trees_din <= x"ffca1615";
		wait for Clk_period;
		Addr <=  "00010101101010";
		Trees_din <= x"008d1615";
		wait for Clk_period;
		Addr <=  "00010101101011";
		Trees_din <= x"ff8d1615";
		wait for Clk_period;
		Addr <=  "00010101101100";
		Trees_din <= x"16000c08";
		wait for Clk_period;
		Addr <=  "00010101101101";
		Trees_din <= x"19008904";
		wait for Clk_period;
		Addr <=  "00010101101110";
		Trees_din <= x"00771615";
		wait for Clk_period;
		Addr <=  "00010101101111";
		Trees_din <= x"ffbc1615";
		wait for Clk_period;
		Addr <=  "00010101110000";
		Trees_din <= x"1702a804";
		wait for Clk_period;
		Addr <=  "00010101110001";
		Trees_din <= x"ff5f1615";
		wait for Clk_period;
		Addr <=  "00010101110010";
		Trees_din <= x"00451615";
		wait for Clk_period;
		Addr <=  "00010101110011";
		Trees_din <= x"20040008";
		wait for Clk_period;
		Addr <=  "00010101110100";
		Trees_din <= x"0200f004";
		wait for Clk_period;
		Addr <=  "00010101110101";
		Trees_din <= x"00ca1615";
		wait for Clk_period;
		Addr <=  "00010101110110";
		Trees_din <= x"00091615";
		wait for Clk_period;
		Addr <=  "00010101110111";
		Trees_din <= x"12fc6f08";
		wait for Clk_period;
		Addr <=  "00010101111000";
		Trees_din <= x"0400ad04";
		wait for Clk_period;
		Addr <=  "00010101111001";
		Trees_din <= x"ff651615";
		wait for Clk_period;
		Addr <=  "00010101111010";
		Trees_din <= x"00371615";
		wait for Clk_period;
		Addr <=  "00010101111011";
		Trees_din <= x"0f00c304";
		wait for Clk_period;
		Addr <=  "00010101111100";
		Trees_din <= x"fffa1615";
		wait for Clk_period;
		Addr <=  "00010101111101";
		Trees_din <= x"001c1615";
		wait for Clk_period;
		Addr <=  "00010101111110";
		Trees_din <= x"0b046008";
		wait for Clk_period;
		Addr <=  "00010101111111";
		Trees_din <= x"10fa6104";
		wait for Clk_period;
		Addr <=  "00010110000000";
		Trees_din <= x"00121615";
		wait for Clk_period;
		Addr <=  "00010110000001";
		Trees_din <= x"007e1615";
		wait for Clk_period;
		Addr <=  "00010110000010";
		Trees_din <= x"000dd204";
		wait for Clk_period;
		Addr <=  "00010110000011";
		Trees_din <= x"00521615";
		wait for Clk_period;
		Addr <=  "00010110000100";
		Trees_din <= x"ffd81615";
		wait for Clk_period;
		Addr <=  "00010110000101";
		Trees_din <= x"01fe6a04";
		wait for Clk_period;
		Addr <=  "00010110000110";
		Trees_din <= x"ff7b16f9";
		wait for Clk_period;
		Addr <=  "00010110000111";
		Trees_din <= x"010d4f34";
		wait for Clk_period;
		Addr <=  "00010110001000";
		Trees_din <= x"03f6f41c";
		wait for Clk_period;
		Addr <=  "00010110001001";
		Trees_din <= x"10028710";
		wait for Clk_period;
		Addr <=  "00010110001010";
		Trees_din <= x"14017208";
		wait for Clk_period;
		Addr <=  "00010110001011";
		Trees_din <= x"1e005b04";
		wait for Clk_period;
		Addr <=  "00010110001100";
		Trees_din <= x"fff416f9";
		wait for Clk_period;
		Addr <=  "00010110001101";
		Trees_din <= x"ff8916f9";
		wait for Clk_period;
		Addr <=  "00010110001110";
		Trees_din <= x"1700f604";
		wait for Clk_period;
		Addr <=  "00010110001111";
		Trees_din <= x"ffff16f9";
		wait for Clk_period;
		Addr <=  "00010110010000";
		Trees_din <= x"013816f9";
		wait for Clk_period;
		Addr <=  "00010110010001";
		Trees_din <= x"04f58908";
		wait for Clk_period;
		Addr <=  "00010110010010";
		Trees_din <= x"16009f04";
		wait for Clk_period;
		Addr <=  "00010110010011";
		Trees_din <= x"000816f9";
		wait for Clk_period;
		Addr <=  "00010110010100";
		Trees_din <= x"ff9b16f9";
		wait for Clk_period;
		Addr <=  "00010110010101";
		Trees_din <= x"ff6216f9";
		wait for Clk_period;
		Addr <=  "00010110010110";
		Trees_din <= x"010d2810";
		wait for Clk_period;
		Addr <=  "00010110010111";
		Trees_din <= x"010cb408";
		wait for Clk_period;
		Addr <=  "00010110011000";
		Trees_din <= x"1703f804";
		wait for Clk_period;
		Addr <=  "00010110011001";
		Trees_din <= x"000216f9";
		wait for Clk_period;
		Addr <=  "00010110011010";
		Trees_din <= x"008316f9";
		wait for Clk_period;
		Addr <=  "00010110011011";
		Trees_din <= x"09005204";
		wait for Clk_period;
		Addr <=  "00010110011100";
		Trees_din <= x"00d616f9";
		wait for Clk_period;
		Addr <=  "00010110011101";
		Trees_din <= x"000e16f9";
		wait for Clk_period;
		Addr <=  "00010110011110";
		Trees_din <= x"02040904";
		wait for Clk_period;
		Addr <=  "00010110011111";
		Trees_din <= x"ff5116f9";
		wait for Clk_period;
		Addr <=  "00010110100000";
		Trees_din <= x"ffd316f9";
		wait for Clk_period;
		Addr <=  "00010110100001";
		Trees_din <= x"03f9d620";
		wait for Clk_period;
		Addr <=  "00010110100010";
		Trees_din <= x"1403ab10";
		wait for Clk_period;
		Addr <=  "00010110100011";
		Trees_din <= x"0f02d608";
		wait for Clk_period;
		Addr <=  "00010110100100";
		Trees_din <= x"08000c04";
		wait for Clk_period;
		Addr <=  "00010110100101";
		Trees_din <= x"ffa716f9";
		wait for Clk_period;
		Addr <=  "00010110100110";
		Trees_din <= x"001616f9";
		wait for Clk_period;
		Addr <=  "00010110100111";
		Trees_din <= x"12027d04";
		wait for Clk_period;
		Addr <=  "00010110101000";
		Trees_din <= x"002016f9";
		wait for Clk_period;
		Addr <=  "00010110101001";
		Trees_din <= x"ff3716f9";
		wait for Clk_period;
		Addr <=  "00010110101010";
		Trees_din <= x"10fade08";
		wait for Clk_period;
		Addr <=  "00010110101011";
		Trees_din <= x"0111ec04";
		wait for Clk_period;
		Addr <=  "00010110101100";
		Trees_din <= x"ff6a16f9";
		wait for Clk_period;
		Addr <=  "00010110101101";
		Trees_din <= x"003e16f9";
		wait for Clk_period;
		Addr <=  "00010110101110";
		Trees_din <= x"0b053004";
		wait for Clk_period;
		Addr <=  "00010110101111";
		Trees_din <= x"00a816f9";
		wait for Clk_period;
		Addr <=  "00010110110000";
		Trees_din <= x"ff9f16f9";
		wait for Clk_period;
		Addr <=  "00010110110001";
		Trees_din <= x"0ef9ce0c";
		wait for Clk_period;
		Addr <=  "00010110110010";
		Trees_din <= x"04fea408";
		wait for Clk_period;
		Addr <=  "00010110110011";
		Trees_din <= x"0a028704";
		wait for Clk_period;
		Addr <=  "00010110110100";
		Trees_din <= x"ffc116f9";
		wait for Clk_period;
		Addr <=  "00010110110101";
		Trees_din <= x"ff1a16f9";
		wait for Clk_period;
		Addr <=  "00010110110110";
		Trees_din <= x"005f16f9";
		wait for Clk_period;
		Addr <=  "00010110110111";
		Trees_din <= x"15008008";
		wait for Clk_period;
		Addr <=  "00010110111000";
		Trees_din <= x"0afcb704";
		wait for Clk_period;
		Addr <=  "00010110111001";
		Trees_din <= x"003d16f9";
		wait for Clk_period;
		Addr <=  "00010110111010";
		Trees_din <= x"ff5716f9";
		wait for Clk_period;
		Addr <=  "00010110111011";
		Trees_din <= x"1400f704";
		wait for Clk_period;
		Addr <=  "00010110111100";
		Trees_din <= x"002316f9";
		wait for Clk_period;
		Addr <=  "00010110111101";
		Trees_din <= x"009316f9";
		wait for Clk_period;
		Addr <=  "00010110111110";
		Trees_din <= x"01fe6a04";
		wait for Clk_period;
		Addr <=  "00010110111111";
		Trees_din <= x"ff7f17d5";
		wait for Clk_period;
		Addr <=  "00010111000000";
		Trees_din <= x"0700563c";
		wait for Clk_period;
		Addr <=  "00010111000001";
		Trees_din <= x"02032e20";
		wait for Clk_period;
		Addr <=  "00010111000010";
		Trees_din <= x"0b047010";
		wait for Clk_period;
		Addr <=  "00010111000011";
		Trees_din <= x"06f96f08";
		wait for Clk_period;
		Addr <=  "00010111000100";
		Trees_din <= x"02fece04";
		wait for Clk_period;
		Addr <=  "00010111000101";
		Trees_din <= x"ffdc17d5";
		wait for Clk_period;
		Addr <=  "00010111000110";
		Trees_din <= x"005017d5";
		wait for Clk_period;
		Addr <=  "00010111000111";
		Trees_din <= x"1a00e504";
		wait for Clk_period;
		Addr <=  "00010111001000";
		Trees_din <= x"fff817d5";
		wait for Clk_period;
		Addr <=  "00010111001001";
		Trees_din <= x"ff6317d5";
		wait for Clk_period;
		Addr <=  "00010111001010";
		Trees_din <= x"09004d08";
		wait for Clk_period;
		Addr <=  "00010111001011";
		Trees_din <= x"01079604";
		wait for Clk_period;
		Addr <=  "00010111001100";
		Trees_din <= x"ffa517d5";
		wait for Clk_period;
		Addr <=  "00010111001101";
		Trees_din <= x"006417d5";
		wait for Clk_period;
		Addr <=  "00010111001110";
		Trees_din <= x"05fe1004";
		wait for Clk_period;
		Addr <=  "00010111001111";
		Trees_din <= x"ff8317d5";
		wait for Clk_period;
		Addr <=  "00010111010000";
		Trees_din <= x"005c17d5";
		wait for Clk_period;
		Addr <=  "00010111010001";
		Trees_din <= x"0d038810";
		wait for Clk_period;
		Addr <=  "00010111010010";
		Trees_din <= x"010b7608";
		wait for Clk_period;
		Addr <=  "00010111010011";
		Trees_din <= x"06f2f004";
		wait for Clk_period;
		Addr <=  "00010111010100";
		Trees_din <= x"003617d5";
		wait for Clk_period;
		Addr <=  "00010111010101";
		Trees_din <= x"ffa417d5";
		wait for Clk_period;
		Addr <=  "00010111010110";
		Trees_din <= x"0afda204";
		wait for Clk_period;
		Addr <=  "00010111010111";
		Trees_din <= x"003a17d5";
		wait for Clk_period;
		Addr <=  "00010111011000";
		Trees_din <= x"ffe417d5";
		wait for Clk_period;
		Addr <=  "00010111011001";
		Trees_din <= x"0002a804";
		wait for Clk_period;
		Addr <=  "00010111011010";
		Trees_din <= x"001417d5";
		wait for Clk_period;
		Addr <=  "00010111011011";
		Trees_din <= x"15009d04";
		wait for Clk_period;
		Addr <=  "00010111011100";
		Trees_din <= x"ff3f17d5";
		wait for Clk_period;
		Addr <=  "00010111011101";
		Trees_din <= x"fff717d5";
		wait for Clk_period;
		Addr <=  "00010111011110";
		Trees_din <= x"18003814";
		wait for Clk_period;
		Addr <=  "00010111011111";
		Trees_din <= x"000b9b08";
		wait for Clk_period;
		Addr <=  "00010111100000";
		Trees_din <= x"16029404";
		wait for Clk_period;
		Addr <=  "00010111100001";
		Trees_din <= x"010817d5";
		wait for Clk_period;
		Addr <=  "00010111100010";
		Trees_din <= x"004a17d5";
		wait for Clk_period;
		Addr <=  "00010111100011";
		Trees_din <= x"08007b04";
		wait for Clk_period;
		Addr <=  "00010111100100";
		Trees_din <= x"00ac17d5";
		wait for Clk_period;
		Addr <=  "00010111100101";
		Trees_din <= x"14019f04";
		wait for Clk_period;
		Addr <=  "00010111100110";
		Trees_din <= x"ffef17d5";
		wait for Clk_period;
		Addr <=  "00010111100111";
		Trees_din <= x"ff9417d5";
		wait for Clk_period;
		Addr <=  "00010111101000";
		Trees_din <= x"1900a410";
		wait for Clk_period;
		Addr <=  "00010111101001";
		Trees_din <= x"15009908";
		wait for Clk_period;
		Addr <=  "00010111101010";
		Trees_din <= x"1e006804";
		wait for Clk_period;
		Addr <=  "00010111101011";
		Trees_din <= x"00b617d5";
		wait for Clk_period;
		Addr <=  "00010111101100";
		Trees_din <= x"001217d5";
		wait for Clk_period;
		Addr <=  "00010111101101";
		Trees_din <= x"1a00d704";
		wait for Clk_period;
		Addr <=  "00010111101110";
		Trees_din <= x"ffde17d5";
		wait for Clk_period;
		Addr <=  "00010111101111";
		Trees_din <= x"005817d5";
		wait for Clk_period;
		Addr <=  "00010111110000";
		Trees_din <= x"07005704";
		wait for Clk_period;
		Addr <=  "00010111110001";
		Trees_din <= x"008517d5";
		wait for Clk_period;
		Addr <=  "00010111110010";
		Trees_din <= x"01107304";
		wait for Clk_period;
		Addr <=  "00010111110011";
		Trees_din <= x"ff9417d5";
		wait for Clk_period;
		Addr <=  "00010111110100";
		Trees_din <= x"004517d5";
		wait for Clk_period;
		Addr <=  "00010111110101";
		Trees_din <= x"01fe6a04";
		wait for Clk_period;
		Addr <=  "00010111110110";
		Trees_din <= x"ff8218c1";
		wait for Clk_period;
		Addr <=  "00010111110111";
		Trees_din <= x"00fd2534";
		wait for Clk_period;
		Addr <=  "00010111111000";
		Trees_din <= x"0f01c21c";
		wait for Clk_period;
		Addr <=  "00010111111001";
		Trees_din <= x"10fbe010";
		wait for Clk_period;
		Addr <=  "00010111111010";
		Trees_din <= x"1900a308";
		wait for Clk_period;
		Addr <=  "00010111111011";
		Trees_din <= x"05fa0504";
		wait for Clk_period;
		Addr <=  "00010111111100";
		Trees_din <= x"fffd18c1";
		wait for Clk_period;
		Addr <=  "00010111111101";
		Trees_din <= x"ffa518c1";
		wait for Clk_period;
		Addr <=  "00010111111110";
		Trees_din <= x"0e017504";
		wait for Clk_period;
		Addr <=  "00010111111111";
		Trees_din <= x"007618c1";
		wait for Clk_period;
		Addr <=  "00011000000000";
		Trees_din <= x"001618c1";
		wait for Clk_period;
		Addr <=  "00011000000001";
		Trees_din <= x"04fd2004";
		wait for Clk_period;
		Addr <=  "00011000000010";
		Trees_din <= x"000b18c1";
		wait for Clk_period;
		Addr <=  "00011000000011";
		Trees_din <= x"07005a04";
		wait for Clk_period;
		Addr <=  "00011000000100";
		Trees_din <= x"ff5c18c1";
		wait for Clk_period;
		Addr <=  "00011000000101";
		Trees_din <= x"ffdf18c1";
		wait for Clk_period;
		Addr <=  "00011000000110";
		Trees_din <= x"00f8f608";
		wait for Clk_period;
		Addr <=  "00011000000111";
		Trees_din <= x"08009104";
		wait for Clk_period;
		Addr <=  "00011000001000";
		Trees_din <= x"00b718c1";
		wait for Clk_period;
		Addr <=  "00011000001001";
		Trees_din <= x"003618c1";
		wait for Clk_period;
		Addr <=  "00011000001010";
		Trees_din <= x"0f031508";
		wait for Clk_period;
		Addr <=  "00011000001011";
		Trees_din <= x"1d004204";
		wait for Clk_period;
		Addr <=  "00011000001100";
		Trees_din <= x"007018c1";
		wait for Clk_period;
		Addr <=  "00011000001101";
		Trees_din <= x"ffef18c1";
		wait for Clk_period;
		Addr <=  "00011000001110";
		Trees_din <= x"0d001504";
		wait for Clk_period;
		Addr <=  "00011000001111";
		Trees_din <= x"000618c1";
		wait for Clk_period;
		Addr <=  "00011000010000";
		Trees_din <= x"ff8718c1";
		wait for Clk_period;
		Addr <=  "00011000010001";
		Trees_din <= x"10f9b120";
		wait for Clk_period;
		Addr <=  "00011000010010";
		Trees_din <= x"0f01a210";
		wait for Clk_period;
		Addr <=  "00011000010011";
		Trees_din <= x"09005308";
		wait for Clk_period;
		Addr <=  "00011000010100";
		Trees_din <= x"010b7604";
		wait for Clk_period;
		Addr <=  "00011000010101";
		Trees_din <= x"ff9c18c1";
		wait for Clk_period;
		Addr <=  "00011000010110";
		Trees_din <= x"007518c1";
		wait for Clk_period;
		Addr <=  "00011000010111";
		Trees_din <= x"19007f04";
		wait for Clk_period;
		Addr <=  "00011000011000";
		Trees_din <= x"005a18c1";
		wait for Clk_period;
		Addr <=  "00011000011001";
		Trees_din <= x"ff7718c1";
		wait for Clk_period;
		Addr <=  "00011000011010";
		Trees_din <= x"16013908";
		wait for Clk_period;
		Addr <=  "00011000011011";
		Trees_din <= x"07005804";
		wait for Clk_period;
		Addr <=  "00011000011100";
		Trees_din <= x"ff7418c1";
		wait for Clk_period;
		Addr <=  "00011000011101";
		Trees_din <= x"003218c1";
		wait for Clk_period;
		Addr <=  "00011000011110";
		Trees_din <= x"03fb3a04";
		wait for Clk_period;
		Addr <=  "00011000011111";
		Trees_din <= x"001718c1";
		wait for Clk_period;
		Addr <=  "00011000100000";
		Trees_din <= x"00d918c1";
		wait for Clk_period;
		Addr <=  "00011000100001";
		Trees_din <= x"14027c10";
		wait for Clk_period;
		Addr <=  "00011000100010";
		Trees_din <= x"03fb9308";
		wait for Clk_period;
		Addr <=  "00011000100011";
		Trees_din <= x"01065e04";
		wait for Clk_period;
		Addr <=  "00011000100100";
		Trees_din <= x"ff8f18c1";
		wait for Clk_period;
		Addr <=  "00011000100101";
		Trees_din <= x"000c18c1";
		wait for Clk_period;
		Addr <=  "00011000100110";
		Trees_din <= x"14024a04";
		wait for Clk_period;
		Addr <=  "00011000100111";
		Trees_din <= x"003118c1";
		wait for Clk_period;
		Addr <=  "00011000101000";
		Trees_din <= x"00cf18c1";
		wait for Clk_period;
		Addr <=  "00011000101001";
		Trees_din <= x"1403b408";
		wait for Clk_period;
		Addr <=  "00011000101010";
		Trees_din <= x"11028704";
		wait for Clk_period;
		Addr <=  "00011000101011";
		Trees_din <= x"fff518c1";
		wait for Clk_period;
		Addr <=  "00011000101100";
		Trees_din <= x"ff9b18c1";
		wait for Clk_period;
		Addr <=  "00011000101101";
		Trees_din <= x"0d000e04";
		wait for Clk_period;
		Addr <=  "00011000101110";
		Trees_din <= x"ffe318c1";
		wait for Clk_period;
		Addr <=  "00011000101111";
		Trees_din <= x"004918c1";
		wait for Clk_period;
		Addr <=  "00011000110000";
		Trees_din <= x"01fe6a04";
		wait for Clk_period;
		Addr <=  "00011000110001";
		Trees_din <= x"ff86197d";
		wait for Clk_period;
		Addr <=  "00011000110010";
		Trees_din <= x"0113e938";
		wait for Clk_period;
		Addr <=  "00011000110011";
		Trees_din <= x"13fa0b18";
		wait for Clk_period;
		Addr <=  "00011000110100";
		Trees_din <= x"0a012808";
		wait for Clk_period;
		Addr <=  "00011000110101";
		Trees_din <= x"1400b604";
		wait for Clk_period;
		Addr <=  "00011000110110";
		Trees_din <= x"fff8197d";
		wait for Clk_period;
		Addr <=  "00011000110111";
		Trees_din <= x"ff5d197d";
		wait for Clk_period;
		Addr <=  "00011000111000";
		Trees_din <= x"05f8c108";
		wait for Clk_period;
		Addr <=  "00011000111001";
		Trees_din <= x"09005504";
		wait for Clk_period;
		Addr <=  "00011000111010";
		Trees_din <= x"0005197d";
		wait for Clk_period;
		Addr <=  "00011000111011";
		Trees_din <= x"ff52197d";
		wait for Clk_period;
		Addr <=  "00011000111100";
		Trees_din <= x"04fa1604";
		wait for Clk_period;
		Addr <=  "00011000111101";
		Trees_din <= x"0057197d";
		wait for Clk_period;
		Addr <=  "00011000111110";
		Trees_din <= x"fff4197d";
		wait for Clk_period;
		Addr <=  "00011000111111";
		Trees_din <= x"13fd6410";
		wait for Clk_period;
		Addr <=  "00011001000000";
		Trees_din <= x"02049a08";
		wait for Clk_period;
		Addr <=  "00011001000001";
		Trees_din <= x"1500a804";
		wait for Clk_period;
		Addr <=  "00011001000010";
		Trees_din <= x"0028197d";
		wait for Clk_period;
		Addr <=  "00011001000011";
		Trees_din <= x"ff68197d";
		wait for Clk_period;
		Addr <=  "00011001000100";
		Trees_din <= x"05fc6904";
		wait for Clk_period;
		Addr <=  "00011001000101";
		Trees_din <= x"00af197d";
		wait for Clk_period;
		Addr <=  "00011001000110";
		Trees_din <= x"ffca197d";
		wait for Clk_period;
		Addr <=  "00011001000111";
		Trees_din <= x"15009908";
		wait for Clk_period;
		Addr <=  "00011001001000";
		Trees_din <= x"1e006804";
		wait for Clk_period;
		Addr <=  "00011001001001";
		Trees_din <= x"005b197d";
		wait for Clk_period;
		Addr <=  "00011001001010";
		Trees_din <= x"0005197d";
		wait for Clk_period;
		Addr <=  "00011001001011";
		Trees_din <= x"1a00e004";
		wait for Clk_period;
		Addr <=  "00011001001100";
		Trees_din <= x"ffd3197d";
		wait for Clk_period;
		Addr <=  "00011001001101";
		Trees_din <= x"001a197d";
		wait for Clk_period;
		Addr <=  "00011001001110";
		Trees_din <= x"1a00e014";
		wait for Clk_period;
		Addr <=  "00011001001111";
		Trees_din <= x"1d004e08";
		wait for Clk_period;
		Addr <=  "00011001010000";
		Trees_din <= x"03f1ef04";
		wait for Clk_period;
		Addr <=  "00011001010001";
		Trees_din <= x"ffee197d";
		wait for Clk_period;
		Addr <=  "00011001010010";
		Trees_din <= x"0089197d";
		wait for Clk_period;
		Addr <=  "00011001010011";
		Trees_din <= x"06f50208";
		wait for Clk_period;
		Addr <=  "00011001010100";
		Trees_din <= x"09005304";
		wait for Clk_period;
		Addr <=  "00011001010101";
		Trees_din <= x"ff9a197d";
		wait for Clk_period;
		Addr <=  "00011001010110";
		Trees_din <= x"fff4197d";
		wait for Clk_period;
		Addr <=  "00011001010111";
		Trees_din <= x"0074197d";
		wait for Clk_period;
		Addr <=  "00011001011000";
		Trees_din <= x"01159308";
		wait for Clk_period;
		Addr <=  "00011001011001";
		Trees_din <= x"13fd9404";
		wait for Clk_period;
		Addr <=  "00011001011010";
		Trees_din <= x"ff85197d";
		wait for Clk_period;
		Addr <=  "00011001011011";
		Trees_din <= x"ffec197d";
		wait for Clk_period;
		Addr <=  "00011001011100";
		Trees_din <= x"0a01c104";
		wait for Clk_period;
		Addr <=  "00011001011101";
		Trees_din <= x"ffe4197d";
		wait for Clk_period;
		Addr <=  "00011001011110";
		Trees_din <= x"0061197d";
		wait for Clk_period;
		Addr <=  "00011001011111";
		Trees_din <= x"01fe6a04";
		wait for Clk_period;
		Addr <=  "00011001100000";
		Trees_din <= x"ff8a19f9";
		wait for Clk_period;
		Addr <=  "00011001100001";
		Trees_din <= x"1703f82c";
		wait for Clk_period;
		Addr <=  "00011001100010";
		Trees_din <= x"1603f918";
		wait for Clk_period;
		Addr <=  "00011001100011";
		Trees_din <= x"1703e110";
		wait for Clk_period;
		Addr <=  "00011001100100";
		Trees_din <= x"07005608";
		wait for Clk_period;
		Addr <=  "00011001100101";
		Trees_din <= x"1005a904";
		wait for Clk_period;
		Addr <=  "00011001100110";
		Trees_din <= x"fffe19f9";
		wait for Clk_period;
		Addr <=  "00011001100111";
		Trees_din <= x"ffa519f9";
		wait for Clk_period;
		Addr <=  "00011001101000";
		Trees_din <= x"1d003904";
		wait for Clk_period;
		Addr <=  "00011001101001";
		Trees_din <= x"008719f9";
		wait for Clk_period;
		Addr <=  "00011001101010";
		Trees_din <= x"000c19f9";
		wait for Clk_period;
		Addr <=  "00011001101011";
		Trees_din <= x"11011c04";
		wait for Clk_period;
		Addr <=  "00011001101100";
		Trees_din <= x"ffec19f9";
		wait for Clk_period;
		Addr <=  "00011001101101";
		Trees_din <= x"00a919f9";
		wait for Clk_period;
		Addr <=  "00011001101110";
		Trees_din <= x"0a040310";
		wait for Clk_period;
		Addr <=  "00011001101111";
		Trees_din <= x"09004508";
		wait for Clk_period;
		Addr <=  "00011001110000";
		Trees_din <= x"1101dc04";
		wait for Clk_period;
		Addr <=  "00011001110001";
		Trees_din <= x"007219f9";
		wait for Clk_period;
		Addr <=  "00011001110010";
		Trees_din <= x"ffc919f9";
		wait for Clk_period;
		Addr <=  "00011001110011";
		Trees_din <= x"0efe4804";
		wait for Clk_period;
		Addr <=  "00011001110100";
		Trees_din <= x"002119f9";
		wait for Clk_period;
		Addr <=  "00011001110101";
		Trees_din <= x"ff8319f9";
		wait for Clk_period;
		Addr <=  "00011001110110";
		Trees_din <= x"00a719f9";
		wait for Clk_period;
		Addr <=  "00011001110111";
		Trees_din <= x"1c002a04";
		wait for Clk_period;
		Addr <=  "00011001111000";
		Trees_din <= x"ff8619f9";
		wait for Clk_period;
		Addr <=  "00011001111001";
		Trees_din <= x"13f85f04";
		wait for Clk_period;
		Addr <=  "00011001111010";
		Trees_din <= x"fffb19f9";
		wait for Clk_period;
		Addr <=  "00011001111011";
		Trees_din <= x"04fd0d04";
		wait for Clk_period;
		Addr <=  "00011001111100";
		Trees_din <= x"003619f9";
		wait for Clk_period;
		Addr <=  "00011001111101";
		Trees_din <= x"00d019f9";
		wait for Clk_period;
		Addr <=  "00011001111110";
		Trees_din <= x"05fcb24c";
		wait for Clk_period;
		Addr <=  "00011001111111";
		Trees_din <= x"05fc5230";
		wait for Clk_period;
		Addr <=  "00011010000000";
		Trees_din <= x"0c001f10";
		wait for Clk_period;
		Addr <=  "00011010000001";
		Trees_din <= x"0209ea0c";
		wait for Clk_period;
		Addr <=  "00011010000010";
		Trees_din <= x"1a00a704";
		wait for Clk_period;
		Addr <=  "00011010000011";
		Trees_din <= x"00041b15";
		wait for Clk_period;
		Addr <=  "00011010000100";
		Trees_din <= x"0e008804";
		wait for Clk_period;
		Addr <=  "00011010000101";
		Trees_din <= x"00cd1b15";
		wait for Clk_period;
		Addr <=  "00011010000110";
		Trees_din <= x"00271b15";
		wait for Clk_period;
		Addr <=  "00011010000111";
		Trees_din <= x"ffab1b15";
		wait for Clk_period;
		Addr <=  "00011010001000";
		Trees_din <= x"0f02f310";
		wait for Clk_period;
		Addr <=  "00011010001001";
		Trees_din <= x"17000108";
		wait for Clk_period;
		Addr <=  "00011010001010";
		Trees_din <= x"0108a404";
		wait for Clk_period;
		Addr <=  "00011010001011";
		Trees_din <= x"ffde1b15";
		wait for Clk_period;
		Addr <=  "00011010001100";
		Trees_din <= x"00521b15";
		wait for Clk_period;
		Addr <=  "00011010001101";
		Trees_din <= x"0f024804";
		wait for Clk_period;
		Addr <=  "00011010001110";
		Trees_din <= x"fff81b15";
		wait for Clk_period;
		Addr <=  "00011010001111";
		Trees_din <= x"00621b15";
		wait for Clk_period;
		Addr <=  "00011010010000";
		Trees_din <= x"19008708";
		wait for Clk_period;
		Addr <=  "00011010010001";
		Trees_din <= x"1a008d04";
		wait for Clk_period;
		Addr <=  "00011010010010";
		Trees_din <= x"ff801b15";
		wait for Clk_period;
		Addr <=  "00011010010011";
		Trees_din <= x"004f1b15";
		wait for Clk_period;
		Addr <=  "00011010010100";
		Trees_din <= x"12027f04";
		wait for Clk_period;
		Addr <=  "00011010010101";
		Trees_din <= x"fff61b15";
		wait for Clk_period;
		Addr <=  "00011010010110";
		Trees_din <= x"ff991b15";
		wait for Clk_period;
		Addr <=  "00011010010111";
		Trees_din <= x"000d6314";
		wait for Clk_period;
		Addr <=  "00011010011000";
		Trees_din <= x"0802ad0c";
		wait for Clk_period;
		Addr <=  "00011010011001";
		Trees_din <= x"0c036e08";
		wait for Clk_period;
		Addr <=  "00011010011010";
		Trees_din <= x"1603f604";
		wait for Clk_period;
		Addr <=  "00011010011011";
		Trees_din <= x"00af1b15";
		wait for Clk_period;
		Addr <=  "00011010011100";
		Trees_din <= x"ffb01b15";
		wait for Clk_period;
		Addr <=  "00011010011101";
		Trees_din <= x"ff8d1b15";
		wait for Clk_period;
		Addr <=  "00011010011110";
		Trees_din <= x"0002d304";
		wait for Clk_period;
		Addr <=  "00011010011111";
		Trees_din <= x"00541b15";
		wait for Clk_period;
		Addr <=  "00011010100000";
		Trees_din <= x"ff5c1b15";
		wait for Clk_period;
		Addr <=  "00011010100001";
		Trees_din <= x"1e005a04";
		wait for Clk_period;
		Addr <=  "00011010100010";
		Trees_din <= x"00201b15";
		wait for Clk_period;
		Addr <=  "00011010100011";
		Trees_din <= x"ff7a1b15";
		wait for Clk_period;
		Addr <=  "00011010100100";
		Trees_din <= x"1102f62c";
		wait for Clk_period;
		Addr <=  "00011010100101";
		Trees_din <= x"1102781c";
		wait for Clk_period;
		Addr <=  "00011010100110";
		Trees_din <= x"0efdd20c";
		wait for Clk_period;
		Addr <=  "00011010100111";
		Trees_din <= x"05fdae04";
		wait for Clk_period;
		Addr <=  "00011010101000";
		Trees_din <= x"ff9a1b15";
		wait for Clk_period;
		Addr <=  "00011010101001";
		Trees_din <= x"0c009c04";
		wait for Clk_period;
		Addr <=  "00011010101010";
		Trees_din <= x"010b1b15";
		wait for Clk_period;
		Addr <=  "00011010101011";
		Trees_din <= x"00301b15";
		wait for Clk_period;
		Addr <=  "00011010101100";
		Trees_din <= x"09005708";
		wait for Clk_period;
		Addr <=  "00011010101101";
		Trees_din <= x"0c014004";
		wait for Clk_period;
		Addr <=  "00011010101110";
		Trees_din <= x"fff71b15";
		wait for Clk_period;
		Addr <=  "00011010101111";
		Trees_din <= x"ff7e1b15";
		wait for Clk_period;
		Addr <=  "00011010110000";
		Trees_din <= x"08005a04";
		wait for Clk_period;
		Addr <=  "00011010110001";
		Trees_din <= x"ffaa1b15";
		wait for Clk_period;
		Addr <=  "00011010110010";
		Trees_din <= x"005f1b15";
		wait for Clk_period;
		Addr <=  "00011010110011";
		Trees_din <= x"06f23704";
		wait for Clk_period;
		Addr <=  "00011010110100";
		Trees_din <= x"00001b15";
		wait for Clk_period;
		Addr <=  "00011010110101";
		Trees_din <= x"19009b04";
		wait for Clk_period;
		Addr <=  "00011010110110";
		Trees_din <= x"ff5c1b15";
		wait for Clk_period;
		Addr <=  "00011010110111";
		Trees_din <= x"01088e04";
		wait for Clk_period;
		Addr <=  "00011010111000";
		Trees_din <= x"ff911b15";
		wait for Clk_period;
		Addr <=  "00011010111001";
		Trees_din <= x"00231b15";
		wait for Clk_period;
		Addr <=  "00011010111010";
		Trees_din <= x"0bf9ce04";
		wait for Clk_period;
		Addr <=  "00011010111011";
		Trees_din <= x"00d91b15";
		wait for Clk_period;
		Addr <=  "00011010111100";
		Trees_din <= x"01045104";
		wait for Clk_period;
		Addr <=  "00011010111101";
		Trees_din <= x"ff851b15";
		wait for Clk_period;
		Addr <=  "00011010111110";
		Trees_din <= x"0200f008";
		wait for Clk_period;
		Addr <=  "00011010111111";
		Trees_din <= x"1e006c04";
		wait for Clk_period;
		Addr <=  "00011011000000";
		Trees_din <= x"00e11b15";
		wait for Clk_period;
		Addr <=  "00011011000001";
		Trees_din <= x"fff81b15";
		wait for Clk_period;
		Addr <=  "00011011000010";
		Trees_din <= x"01096904";
		wait for Clk_period;
		Addr <=  "00011011000011";
		Trees_din <= x"ff931b15";
		wait for Clk_period;
		Addr <=  "00011011000100";
		Trees_din <= x"00191b15";
		wait for Clk_period;
		Addr <=  "00011011000101";
		Trees_din <= x"20040034";
		wait for Clk_period;
		Addr <=  "00011011000110";
		Trees_din <= x"05f9a418";
		wait for Clk_period;
		Addr <=  "00011011000111";
		Trees_din <= x"19009e14";
		wait for Clk_period;
		Addr <=  "00011011001000";
		Trees_din <= x"0014870c";
		wait for Clk_period;
		Addr <=  "00011011001001";
		Trees_din <= x"02077508";
		wait for Clk_period;
		Addr <=  "00011011001010";
		Trees_din <= x"02ffb904";
		wait for Clk_period;
		Addr <=  "00011011001011";
		Trees_din <= x"ffe31c29";
		wait for Clk_period;
		Addr <=  "00011011001100";
		Trees_din <= x"00b01c29";
		wait for Clk_period;
		Addr <=  "00011011001101";
		Trees_din <= x"ffcd1c29";
		wait for Clk_period;
		Addr <=  "00011011001110";
		Trees_din <= x"0f023404";
		wait for Clk_period;
		Addr <=  "00011011001111";
		Trees_din <= x"00121c29";
		wait for Clk_period;
		Addr <=  "00011011010000";
		Trees_din <= x"ffb61c29";
		wait for Clk_period;
		Addr <=  "00011011010001";
		Trees_din <= x"ffa51c29";
		wait for Clk_period;
		Addr <=  "00011011010010";
		Trees_din <= x"1103d614";
		wait for Clk_period;
		Addr <=  "00011011010011";
		Trees_din <= x"18004f0c";
		wait for Clk_period;
		Addr <=  "00011011010100";
		Trees_din <= x"010fd308";
		wait for Clk_period;
		Addr <=  "00011011010101";
		Trees_din <= x"11ff2e04";
		wait for Clk_period;
		Addr <=  "00011011010110";
		Trees_din <= x"ffdf1c29";
		wait for Clk_period;
		Addr <=  "00011011010111";
		Trees_din <= x"ff4f1c29";
		wait for Clk_period;
		Addr <=  "00011011011000";
		Trees_din <= x"00261c29";
		wait for Clk_period;
		Addr <=  "00011011011001";
		Trees_din <= x"1600b804";
		wait for Clk_period;
		Addr <=  "00011011011010";
		Trees_din <= x"007f1c29";
		wait for Clk_period;
		Addr <=  "00011011011011";
		Trees_din <= x"ff931c29";
		wait for Clk_period;
		Addr <=  "00011011011100";
		Trees_din <= x"02010204";
		wait for Clk_period;
		Addr <=  "00011011011101";
		Trees_din <= x"009a1c29";
		wait for Clk_period;
		Addr <=  "00011011011110";
		Trees_din <= x"ffb11c29";
		wait for Clk_period;
		Addr <=  "00011011011111";
		Trees_din <= x"03f36e20";
		wait for Clk_period;
		Addr <=  "00011011100000";
		Trees_din <= x"1d004a10";
		wait for Clk_period;
		Addr <=  "00011011100001";
		Trees_din <= x"1f00010c";
		wait for Clk_period;
		Addr <=  "00011011100010";
		Trees_din <= x"04f62904";
		wait for Clk_period;
		Addr <=  "00011011100011";
		Trees_din <= x"ff8a1c29";
		wait for Clk_period;
		Addr <=  "00011011100100";
		Trees_din <= x"13fe1b04";
		wait for Clk_period;
		Addr <=  "00011011100101";
		Trees_din <= x"006b1c29";
		wait for Clk_period;
		Addr <=  "00011011100110";
		Trees_din <= x"ffbd1c29";
		wait for Clk_period;
		Addr <=  "00011011100111";
		Trees_din <= x"006d1c29";
		wait for Clk_period;
		Addr <=  "00011011101000";
		Trees_din <= x"03f1ef04";
		wait for Clk_period;
		Addr <=  "00011011101001";
		Trees_din <= x"ffed1c29";
		wait for Clk_period;
		Addr <=  "00011011101010";
		Trees_din <= x"1c003c04";
		wait for Clk_period;
		Addr <=  "00011011101011";
		Trees_din <= x"01341c29";
		wait for Clk_period;
		Addr <=  "00011011101100";
		Trees_din <= x"0a01db04";
		wait for Clk_period;
		Addr <=  "00011011101101";
		Trees_din <= x"00251c29";
		wait for Clk_period;
		Addr <=  "00011011101110";
		Trees_din <= x"00981c29";
		wait for Clk_period;
		Addr <=  "00011011101111";
		Trees_din <= x"1e005b1c";
		wait for Clk_period;
		Addr <=  "00011011110000";
		Trees_din <= x"1201e20c";
		wait for Clk_period;
		Addr <=  "00011011110001";
		Trees_din <= x"15009904";
		wait for Clk_period;
		Addr <=  "00011011110010";
		Trees_din <= x"00b71c29";
		wait for Clk_period;
		Addr <=  "00011011110011";
		Trees_din <= x"08004404";
		wait for Clk_period;
		Addr <=  "00011011110100";
		Trees_din <= x"00611c29";
		wait for Clk_period;
		Addr <=  "00011011110101";
		Trees_din <= x"ffc91c29";
		wait for Clk_period;
		Addr <=  "00011011110110";
		Trees_din <= x"14027c08";
		wait for Clk_period;
		Addr <=  "00011011110111";
		Trees_din <= x"10055404";
		wait for Clk_period;
		Addr <=  "00011011111000";
		Trees_din <= x"007d1c29";
		wait for Clk_period;
		Addr <=  "00011011111001";
		Trees_din <= x"ffd41c29";
		wait for Clk_period;
		Addr <=  "00011011111010";
		Trees_din <= x"05fc0404";
		wait for Clk_period;
		Addr <=  "00011011111011";
		Trees_din <= x"ff9d1c29";
		wait for Clk_period;
		Addr <=  "00011011111100";
		Trees_din <= x"007b1c29";
		wait for Clk_period;
		Addr <=  "00011011111101";
		Trees_din <= x"1800390c";
		wait for Clk_period;
		Addr <=  "00011011111110";
		Trees_din <= x"1b003204";
		wait for Clk_period;
		Addr <=  "00011011111111";
		Trees_din <= x"ff3d1c29";
		wait for Clk_period;
		Addr <=  "00011100000000";
		Trees_din <= x"1b003304";
		wait for Clk_period;
		Addr <=  "00011100000001";
		Trees_din <= x"000d1c29";
		wait for Clk_period;
		Addr <=  "00011100000010";
		Trees_din <= x"ff9d1c29";
		wait for Clk_period;
		Addr <=  "00011100000011";
		Trees_din <= x"1301ab08";
		wait for Clk_period;
		Addr <=  "00011100000100";
		Trees_din <= x"12028604";
		wait for Clk_period;
		Addr <=  "00011100000101";
		Trees_din <= x"00091c29";
		wait for Clk_period;
		Addr <=  "00011100000110";
		Trees_din <= x"ffd21c29";
		wait for Clk_period;
		Addr <=  "00011100000111";
		Trees_din <= x"06f74a04";
		wait for Clk_period;
		Addr <=  "00011100001000";
		Trees_din <= x"007f1c29";
		wait for Clk_period;
		Addr <=  "00011100001001";
		Trees_din <= x"ffb71c29";
		wait for Clk_period;
		Addr <=  "00011100001010";
		Trees_din <= x"01fe6a04";
		wait for Clk_period;
		Addr <=  "00011100001011";
		Trees_din <= x"ff901ced";
		wait for Clk_period;
		Addr <=  "00011100001100";
		Trees_din <= x"0113e93c";
		wait for Clk_period;
		Addr <=  "00011100001101";
		Trees_din <= x"0bf9231c";
		wait for Clk_period;
		Addr <=  "00011100001110";
		Trees_din <= x"09005610";
		wait for Clk_period;
		Addr <=  "00011100001111";
		Trees_din <= x"01090e08";
		wait for Clk_period;
		Addr <=  "00011100010000";
		Trees_din <= x"19009d04";
		wait for Clk_period;
		Addr <=  "00011100010001";
		Trees_din <= x"ffee1ced";
		wait for Clk_period;
		Addr <=  "00011100010010";
		Trees_din <= x"ff891ced";
		wait for Clk_period;
		Addr <=  "00011100010011";
		Trees_din <= x"03f85a04";
		wait for Clk_period;
		Addr <=  "00011100010100";
		Trees_din <= x"fffd1ced";
		wait for Clk_period;
		Addr <=  "00011100010101";
		Trees_din <= x"00941ced";
		wait for Clk_period;
		Addr <=  "00011100010110";
		Trees_din <= x"11013d08";
		wait for Clk_period;
		Addr <=  "00011100010111";
		Trees_din <= x"0c02cf04";
		wait for Clk_period;
		Addr <=  "00011100011000";
		Trees_din <= x"003e1ced";
		wait for Clk_period;
		Addr <=  "00011100011001";
		Trees_din <= x"ffc71ced";
		wait for Clk_period;
		Addr <=  "00011100011010";
		Trees_din <= x"ff511ced";
		wait for Clk_period;
		Addr <=  "00011100011011";
		Trees_din <= x"1500a010";
		wait for Clk_period;
		Addr <=  "00011100011100";
		Trees_din <= x"18003c08";
		wait for Clk_period;
		Addr <=  "00011100011101";
		Trees_din <= x"0afaf204";
		wait for Clk_period;
		Addr <=  "00011100011110";
		Trees_din <= x"ffbf1ced";
		wait for Clk_period;
		Addr <=  "00011100011111";
		Trees_din <= x"006f1ced";
		wait for Clk_period;
		Addr <=  "00011100100000";
		Trees_din <= x"13025704";
		wait for Clk_period;
		Addr <=  "00011100100001";
		Trees_din <= x"00021ced";
		wait for Clk_period;
		Addr <=  "00011100100010";
		Trees_din <= x"00571ced";
		wait for Clk_period;
		Addr <=  "00011100100011";
		Trees_din <= x"1500a408";
		wait for Clk_period;
		Addr <=  "00011100100100";
		Trees_din <= x"1c003104";
		wait for Clk_period;
		Addr <=  "00011100100101";
		Trees_din <= x"ff8a1ced";
		wait for Clk_period;
		Addr <=  "00011100100110";
		Trees_din <= x"002c1ced";
		wait for Clk_period;
		Addr <=  "00011100100111";
		Trees_din <= x"11045b04";
		wait for Clk_period;
		Addr <=  "00011100101000";
		Trees_din <= x"fffe1ced";
		wait for Clk_period;
		Addr <=  "00011100101001";
		Trees_din <= x"00951ced";
		wait for Clk_period;
		Addr <=  "00011100101010";
		Trees_din <= x"1a00e014";
		wait for Clk_period;
		Addr <=  "00011100101011";
		Trees_din <= x"1d004f08";
		wait for Clk_period;
		Addr <=  "00011100101100";
		Trees_din <= x"0015f004";
		wait for Clk_period;
		Addr <=  "00011100101101";
		Trees_din <= x"00881ced";
		wait for Clk_period;
		Addr <=  "00011100101110";
		Trees_din <= x"000a1ced";
		wait for Clk_period;
		Addr <=  "00011100101111";
		Trees_din <= x"06f50208";
		wait for Clk_period;
		Addr <=  "00011100110000";
		Trees_din <= x"09005304";
		wait for Clk_period;
		Addr <=  "00011100110001";
		Trees_din <= x"ffa11ced";
		wait for Clk_period;
		Addr <=  "00011100110010";
		Trees_din <= x"fff41ced";
		wait for Clk_period;
		Addr <=  "00011100110011";
		Trees_din <= x"00691ced";
		wait for Clk_period;
		Addr <=  "00011100110100";
		Trees_din <= x"01159308";
		wait for Clk_period;
		Addr <=  "00011100110101";
		Trees_din <= x"0a026704";
		wait for Clk_period;
		Addr <=  "00011100110110";
		Trees_din <= x"ffec1ced";
		wait for Clk_period;
		Addr <=  "00011100110111";
		Trees_din <= x"ff991ced";
		wait for Clk_period;
		Addr <=  "00011100111000";
		Trees_din <= x"0a023504";
		wait for Clk_period;
		Addr <=  "00011100111001";
		Trees_din <= x"ffec1ced";
		wait for Clk_period;
		Addr <=  "00011100111010";
		Trees_din <= x"005a1ced";
		wait for Clk_period;
		Addr <=  "00011100111011";
		Trees_din <= x"0c03cc68";
		wait for Clk_period;
		Addr <=  "00011100111100";
		Trees_din <= x"010f7440";
		wait for Clk_period;
		Addr <=  "00011100111101";
		Trees_din <= x"0f005020";
		wait for Clk_period;
		Addr <=  "00011100111110";
		Trees_din <= x"17000810";
		wait for Clk_period;
		Addr <=  "00011100111111";
		Trees_din <= x"04faa908";
		wait for Clk_period;
		Addr <=  "00011101000000";
		Trees_din <= x"13ff6104";
		wait for Clk_period;
		Addr <=  "00011101000001";
		Trees_din <= x"00031e09";
		wait for Clk_period;
		Addr <=  "00011101000010";
		Trees_din <= x"00e11e09";
		wait for Clk_period;
		Addr <=  "00011101000011";
		Trees_din <= x"12028204";
		wait for Clk_period;
		Addr <=  "00011101000100";
		Trees_din <= x"ff8e1e09";
		wait for Clk_period;
		Addr <=  "00011101000101";
		Trees_din <= x"00751e09";
		wait for Clk_period;
		Addr <=  "00011101000110";
		Trees_din <= x"0e037808";
		wait for Clk_period;
		Addr <=  "00011101000111";
		Trees_din <= x"17006004";
		wait for Clk_period;
		Addr <=  "00011101001000";
		Trees_din <= x"ff7f1e09";
		wait for Clk_period;
		Addr <=  "00011101001001";
		Trees_din <= x"fff41e09";
		wait for Clk_period;
		Addr <=  "00011101001010";
		Trees_din <= x"07005a04";
		wait for Clk_period;
		Addr <=  "00011101001011";
		Trees_din <= x"ff4f1e09";
		wait for Clk_period;
		Addr <=  "00011101001100";
		Trees_din <= x"ffd81e09";
		wait for Clk_period;
		Addr <=  "00011101001101";
		Trees_din <= x"14027c10";
		wait for Clk_period;
		Addr <=  "00011101001110";
		Trees_din <= x"1c003d08";
		wait for Clk_period;
		Addr <=  "00011101001111";
		Trees_din <= x"1900a704";
		wait for Clk_period;
		Addr <=  "00011101010000";
		Trees_din <= x"00401e09";
		wait for Clk_period;
		Addr <=  "00011101010001";
		Trees_din <= x"ffdc1e09";
		wait for Clk_period;
		Addr <=  "00011101010010";
		Trees_din <= x"02039104";
		wait for Clk_period;
		Addr <=  "00011101010011";
		Trees_din <= x"000f1e09";
		wait for Clk_period;
		Addr <=  "00011101010100";
		Trees_din <= x"ff991e09";
		wait for Clk_period;
		Addr <=  "00011101010101";
		Trees_din <= x"1403b408";
		wait for Clk_period;
		Addr <=  "00011101010110";
		Trees_din <= x"0407e104";
		wait for Clk_period;
		Addr <=  "00011101010111";
		Trees_din <= x"ffb51e09";
		wait for Clk_period;
		Addr <=  "00011101011000";
		Trees_din <= x"003a1e09";
		wait for Clk_period;
		Addr <=  "00011101011001";
		Trees_din <= x"0d001204";
		wait for Clk_period;
		Addr <=  "00011101011010";
		Trees_din <= x"ffd31e09";
		wait for Clk_period;
		Addr <=  "00011101011011";
		Trees_din <= x"00411e09";
		wait for Clk_period;
		Addr <=  "00011101011100";
		Trees_din <= x"07005c1c";
		wait for Clk_period;
		Addr <=  "00011101011101";
		Trees_din <= x"03f9f210";
		wait for Clk_period;
		Addr <=  "00011101011110";
		Trees_din <= x"0a02f108";
		wait for Clk_period;
		Addr <=  "00011101011111";
		Trees_din <= x"0c00aa04";
		wait for Clk_period;
		Addr <=  "00011101100000";
		Trees_din <= x"00581e09";
		wait for Clk_period;
		Addr <=  "00011101100001";
		Trees_din <= x"fff51e09";
		wait for Clk_period;
		Addr <=  "00011101100010";
		Trees_din <= x"04f72f04";
		wait for Clk_period;
		Addr <=  "00011101100011";
		Trees_din <= x"00661e09";
		wait for Clk_period;
		Addr <=  "00011101100100";
		Trees_din <= x"ff7f1e09";
		wait for Clk_period;
		Addr <=  "00011101100101";
		Trees_din <= x"0ef9ce04";
		wait for Clk_period;
		Addr <=  "00011101100110";
		Trees_din <= x"ffd51e09";
		wait for Clk_period;
		Addr <=  "00011101100111";
		Trees_din <= x"00005104";
		wait for Clk_period;
		Addr <=  "00011101101000";
		Trees_din <= x"000a1e09";
		wait for Clk_period;
		Addr <=  "00011101101001";
		Trees_din <= x"008f1e09";
		wait for Clk_period;
		Addr <=  "00011101101010";
		Trees_din <= x"04f73904";
		wait for Clk_period;
		Addr <=  "00011101101011";
		Trees_din <= x"fffc1e09";
		wait for Clk_period;
		Addr <=  "00011101101100";
		Trees_din <= x"1e007e04";
		wait for Clk_period;
		Addr <=  "00011101101101";
		Trees_din <= x"00ae1e09";
		wait for Clk_period;
		Addr <=  "00011101101110";
		Trees_din <= x"00311e09";
		wait for Clk_period;
		Addr <=  "00011101101111";
		Trees_din <= x"0d013608";
		wait for Clk_period;
		Addr <=  "00011101110000";
		Trees_din <= x"03f97304";
		wait for Clk_period;
		Addr <=  "00011101110001";
		Trees_din <= x"000f1e09";
		wait for Clk_period;
		Addr <=  "00011101110010";
		Trees_din <= x"ff881e09";
		wait for Clk_period;
		Addr <=  "00011101110011";
		Trees_din <= x"12005e0c";
		wait for Clk_period;
		Addr <=  "00011101110100";
		Trees_din <= x"0209bd08";
		wait for Clk_period;
		Addr <=  "00011101110101";
		Trees_din <= x"02058f04";
		wait for Clk_period;
		Addr <=  "00011101110110";
		Trees_din <= x"ffec1e09";
		wait for Clk_period;
		Addr <=  "00011101110111";
		Trees_din <= x"ff681e09";
		wait for Clk_period;
		Addr <=  "00011101111000";
		Trees_din <= x"00561e09";
		wait for Clk_period;
		Addr <=  "00011101111001";
		Trees_din <= x"0c03ee08";
		wait for Clk_period;
		Addr <=  "00011101111010";
		Trees_din <= x"15009d04";
		wait for Clk_period;
		Addr <=  "00011101111011";
		Trees_din <= x"00cd1e09";
		wait for Clk_period;
		Addr <=  "00011101111100";
		Trees_din <= x"002c1e09";
		wait for Clk_period;
		Addr <=  "00011101111101";
		Trees_din <= x"03f9b804";
		wait for Clk_period;
		Addr <=  "00011101111110";
		Trees_din <= x"ffa51e09";
		wait for Clk_period;
		Addr <=  "00011101111111";
		Trees_din <= x"01067004";
		wait for Clk_period;
		Addr <=  "00011110000000";
		Trees_din <= x"00061e09";
		wait for Clk_period;
		Addr <=  "00011110000001";
		Trees_din <= x"006e1e09";
		wait for Clk_period;
		Addr <=  "00011110000010";
		Trees_din <= x"1a00810c";
		wait for Clk_period;
		Addr <=  "00011110000011";
		Trees_din <= x"03f91104";
		wait for Clk_period;
		Addr <=  "00011110000100";
		Trees_din <= x"ffdb1e7d";
		wait for Clk_period;
		Addr <=  "00011110000101";
		Trees_din <= x"04f9f304";
		wait for Clk_period;
		Addr <=  "00011110000110";
		Trees_din <= x"00b91e7d";
		wait for Clk_period;
		Addr <=  "00011110000111";
		Trees_din <= x"00151e7d";
		wait for Clk_period;
		Addr <=  "00011110001000";
		Trees_din <= x"18005528";
		wait for Clk_period;
		Addr <=  "00011110001001";
		Trees_din <= x"1d005820";
		wait for Clk_period;
		Addr <=  "00011110001010";
		Trees_din <= x"0d03bf10";
		wait for Clk_period;
		Addr <=  "00011110001011";
		Trees_din <= x"0d02c808";
		wait for Clk_period;
		Addr <=  "00011110001100";
		Trees_din <= x"0d021904";
		wait for Clk_period;
		Addr <=  "00011110001101";
		Trees_din <= x"00091e7d";
		wait for Clk_period;
		Addr <=  "00011110001110";
		Trees_din <= x"ffc71e7d";
		wait for Clk_period;
		Addr <=  "00011110001111";
		Trees_din <= x"0b057c04";
		wait for Clk_period;
		Addr <=  "00011110010000";
		Trees_din <= x"000d1e7d";
		wait for Clk_period;
		Addr <=  "00011110010001";
		Trees_din <= x"00af1e7d";
		wait for Clk_period;
		Addr <=  "00011110010010";
		Trees_din <= x"07005908";
		wait for Clk_period;
		Addr <=  "00011110010011";
		Trees_din <= x"0200e804";
		wait for Clk_period;
		Addr <=  "00011110010100";
		Trees_din <= x"00091e7d";
		wait for Clk_period;
		Addr <=  "00011110010101";
		Trees_din <= x"ff6c1e7d";
		wait for Clk_period;
		Addr <=  "00011110010110";
		Trees_din <= x"00054504";
		wait for Clk_period;
		Addr <=  "00011110010111";
		Trees_din <= x"ffc01e7d";
		wait for Clk_period;
		Addr <=  "00011110011000";
		Trees_din <= x"00511e7d";
		wait for Clk_period;
		Addr <=  "00011110011001";
		Trees_din <= x"010c6804";
		wait for Clk_period;
		Addr <=  "00011110011010";
		Trees_din <= x"ffeb1e7d";
		wait for Clk_period;
		Addr <=  "00011110011011";
		Trees_din <= x"00b01e7d";
		wait for Clk_period;
		Addr <=  "00011110011100";
		Trees_din <= x"08002604";
		wait for Clk_period;
		Addr <=  "00011110011101";
		Trees_din <= x"fffb1e7d";
		wait for Clk_period;
		Addr <=  "00011110011110";
		Trees_din <= x"ff681e7d";
		wait for Clk_period;
		Addr <=  "00011110011111";
		Trees_din <= x"0118034c";
		wait for Clk_period;
		Addr <=  "00011110100000";
		Trees_din <= x"10f72510";
		wait for Clk_period;
		Addr <=  "00011110100001";
		Trees_din <= x"00042108";
		wait for Clk_period;
		Addr <=  "00011110100010";
		Trees_din <= x"0a02ad04";
		wait for Clk_period;
		Addr <=  "00011110100011";
		Trees_din <= x"001e1f19";
		wait for Clk_period;
		Addr <=  "00011110100100";
		Trees_din <= x"00b01f19";
		wait for Clk_period;
		Addr <=  "00011110100101";
		Trees_din <= x"010d9004";
		wait for Clk_period;
		Addr <=  "00011110100110";
		Trees_din <= x"ff851f19";
		wait for Clk_period;
		Addr <=  "00011110100111";
		Trees_din <= x"00701f19";
		wait for Clk_period;
		Addr <=  "00011110101000";
		Trees_din <= x"10f9b11c";
		wait for Clk_period;
		Addr <=  "00011110101001";
		Trees_din <= x"05f8c10c";
		wait for Clk_period;
		Addr <=  "00011110101010";
		Trees_din <= x"0011cf08";
		wait for Clk_period;
		Addr <=  "00011110101011";
		Trees_din <= x"1d004104";
		wait for Clk_period;
		Addr <=  "00011110101100";
		Trees_din <= x"000d1f19";
		wait for Clk_period;
		Addr <=  "00011110101101";
		Trees_din <= x"00aa1f19";
		wait for Clk_period;
		Addr <=  "00011110101110";
		Trees_din <= x"ffe01f19";
		wait for Clk_period;
		Addr <=  "00011110101111";
		Trees_din <= x"03f71408";
		wait for Clk_period;
		Addr <=  "00011110110000";
		Trees_din <= x"04f9f304";
		wait for Clk_period;
		Addr <=  "00011110110001";
		Trees_din <= x"ffba1f19";
		wait for Clk_period;
		Addr <=  "00011110110010";
		Trees_din <= x"00b61f19";
		wait for Clk_period;
		Addr <=  "00011110110011";
		Trees_din <= x"0f01af04";
		wait for Clk_period;
		Addr <=  "00011110110100";
		Trees_din <= x"ff861f19";
		wait for Clk_period;
		Addr <=  "00011110110101";
		Trees_din <= x"fffa1f19";
		wait for Clk_period;
		Addr <=  "00011110110110";
		Trees_din <= x"10fa3b10";
		wait for Clk_period;
		Addr <=  "00011110110111";
		Trees_din <= x"16009f08";
		wait for Clk_period;
		Addr <=  "00011110111000";
		Trees_din <= x"0afcf304";
		wait for Clk_period;
		Addr <=  "00011110111001";
		Trees_din <= x"007e1f19";
		wait for Clk_period;
		Addr <=  "00011110111010";
		Trees_din <= x"ff751f19";
		wait for Clk_period;
		Addr <=  "00011110111011";
		Trees_din <= x"1402e804";
		wait for Clk_period;
		Addr <=  "00011110111100";
		Trees_din <= x"008b1f19";
		wait for Clk_period;
		Addr <=  "00011110111101";
		Trees_din <= x"ffd31f19";
		wait for Clk_period;
		Addr <=  "00011110111110";
		Trees_din <= x"0302da08";
		wait for Clk_period;
		Addr <=  "00011110111111";
		Trees_din <= x"09005b04";
		wait for Clk_period;
		Addr <=  "00011111000000";
		Trees_din <= x"00091f19";
		wait for Clk_period;
		Addr <=  "00011111000001";
		Trees_din <= x"ffc91f19";
		wait for Clk_period;
		Addr <=  "00011111000010";
		Trees_din <= x"04f83e04";
		wait for Clk_period;
		Addr <=  "00011111000011";
		Trees_din <= x"00681f19";
		wait for Clk_period;
		Addr <=  "00011111000100";
		Trees_din <= x"ffba1f19";
		wait for Clk_period;
		Addr <=  "00011111000101";
		Trees_din <= x"006c1f19";
		wait for Clk_period;
		Addr <=  "00011111000110";
		Trees_din <= x"15009930";
		wait for Clk_period;
		Addr <=  "00011111000111";
		Trees_din <= x"18003d0c";
		wait for Clk_period;
		Addr <=  "00011111001000";
		Trees_din <= x"1900a404";
		wait for Clk_period;
		Addr <=  "00011111001001";
		Trees_din <= x"00d82035";
		wait for Clk_period;
		Addr <=  "00011111001010";
		Trees_din <= x"1900b404";
		wait for Clk_period;
		Addr <=  "00011111001011";
		Trees_din <= x"ffd82035";
		wait for Clk_period;
		Addr <=  "00011111001100";
		Trees_din <= x"00512035";
		wait for Clk_period;
		Addr <=  "00011111001101";
		Trees_din <= x"1900aa20";
		wait for Clk_period;
		Addr <=  "00011111001110";
		Trees_din <= x"15009010";
		wait for Clk_period;
		Addr <=  "00011111001111";
		Trees_din <= x"0d030d08";
		wait for Clk_period;
		Addr <=  "00011111010000";
		Trees_din <= x"010f0b04";
		wait for Clk_period;
		Addr <=  "00011111010001";
		Trees_din <= x"fff82035";
		wait for Clk_period;
		Addr <=  "00011111010010";
		Trees_din <= x"00452035";
		wait for Clk_period;
		Addr <=  "00011111010011";
		Trees_din <= x"1c003f04";
		wait for Clk_period;
		Addr <=  "00011111010100";
		Trees_din <= x"ff892035";
		wait for Clk_period;
		Addr <=  "00011111010101";
		Trees_din <= x"00042035";
		wait for Clk_period;
		Addr <=  "00011111010110";
		Trees_din <= x"0c00db08";
		wait for Clk_period;
		Addr <=  "00011111010111";
		Trees_din <= x"08007b04";
		wait for Clk_period;
		Addr <=  "00011111011000";
		Trees_din <= x"001f2035";
		wait for Clk_period;
		Addr <=  "00011111011001";
		Trees_din <= x"ff982035";
		wait for Clk_period;
		Addr <=  "00011111011010";
		Trees_din <= x"0103f604";
		wait for Clk_period;
		Addr <=  "00011111011011";
		Trees_din <= x"ffa42035";
		wait for Clk_period;
		Addr <=  "00011111011100";
		Trees_din <= x"00452035";
		wait for Clk_period;
		Addr <=  "00011111011101";
		Trees_din <= x"ff6f2035";
		wait for Clk_period;
		Addr <=  "00011111011110";
		Trees_din <= x"0111ec40";
		wait for Clk_period;
		Addr <=  "00011111011111";
		Trees_din <= x"1e006420";
		wait for Clk_period;
		Addr <=  "00011111100000";
		Trees_din <= x"1201e210";
		wait for Clk_period;
		Addr <=  "00011111100001";
		Trees_din <= x"07005608";
		wait for Clk_period;
		Addr <=  "00011111100010";
		Trees_din <= x"02fcb504";
		wait for Clk_period;
		Addr <=  "00011111100011";
		Trees_din <= x"00502035";
		wait for Clk_period;
		Addr <=  "00011111100100";
		Trees_din <= x"ffb42035";
		wait for Clk_period;
		Addr <=  "00011111100101";
		Trees_din <= x"03011204";
		wait for Clk_period;
		Addr <=  "00011111100110";
		Trees_din <= x"002d2035";
		wait for Clk_period;
		Addr <=  "00011111100111";
		Trees_din <= x"ffaf2035";
		wait for Clk_period;
		Addr <=  "00011111101000";
		Trees_din <= x"11048708";
		wait for Clk_period;
		Addr <=  "00011111101001";
		Trees_din <= x"06f1d904";
		wait for Clk_period;
		Addr <=  "00011111101010";
		Trees_din <= x"008a2035";
		wait for Clk_period;
		Addr <=  "00011111101011";
		Trees_din <= x"00032035";
		wait for Clk_period;
		Addr <=  "00011111101100";
		Trees_din <= x"18003b04";
		wait for Clk_period;
		Addr <=  "00011111101101";
		Trees_din <= x"00b52035";
		wait for Clk_period;
		Addr <=  "00011111101110";
		Trees_din <= x"00262035";
		wait for Clk_period;
		Addr <=  "00011111101111";
		Trees_din <= x"1e006a10";
		wait for Clk_period;
		Addr <=  "00011111110000";
		Trees_din <= x"0bf92c08";
		wait for Clk_period;
		Addr <=  "00011111110001";
		Trees_din <= x"0800f004";
		wait for Clk_period;
		Addr <=  "00011111110010";
		Trees_din <= x"ffde2035";
		wait for Clk_period;
		Addr <=  "00011111110011";
		Trees_din <= x"00822035";
		wait for Clk_period;
		Addr <=  "00011111110100";
		Trees_din <= x"05fc4404";
		wait for Clk_period;
		Addr <=  "00011111110101";
		Trees_din <= x"ff712035";
		wait for Clk_period;
		Addr <=  "00011111110110";
		Trees_din <= x"ffef2035";
		wait for Clk_period;
		Addr <=  "00011111110111";
		Trees_din <= x"11029208";
		wait for Clk_period;
		Addr <=  "00011111111000";
		Trees_din <= x"04fe8104";
		wait for Clk_period;
		Addr <=  "00011111111001";
		Trees_din <= x"00612035";
		wait for Clk_period;
		Addr <=  "00011111111010";
		Trees_din <= x"ffc72035";
		wait for Clk_period;
		Addr <=  "00011111111011";
		Trees_din <= x"03fc2f04";
		wait for Clk_period;
		Addr <=  "00011111111100";
		Trees_din <= x"ff7b2035";
		wait for Clk_period;
		Addr <=  "00011111111101";
		Trees_din <= x"00392035";
		wait for Clk_period;
		Addr <=  "00011111111110";
		Trees_din <= x"05f7e710";
		wait for Clk_period;
		Addr <=  "00011111111111";
		Trees_din <= x"000b9b04";
		wait for Clk_period;
		Addr <=  "00100000000000";
		Trees_din <= x"005e2035";
		wait for Clk_period;
		Addr <=  "00100000000001";
		Trees_din <= x"01159308";
		wait for Clk_period;
		Addr <=  "00100000000010";
		Trees_din <= x"0e008204";
		wait for Clk_period;
		Addr <=  "00100000000011";
		Trees_din <= x"ff7d2035";
		wait for Clk_period;
		Addr <=  "00100000000100";
		Trees_din <= x"ffdf2035";
		wait for Clk_period;
		Addr <=  "00100000000101";
		Trees_din <= x"00242035";
		wait for Clk_period;
		Addr <=  "00100000000110";
		Trees_din <= x"09005708";
		wait for Clk_period;
		Addr <=  "00100000000111";
		Trees_din <= x"01123c04";
		wait for Clk_period;
		Addr <=  "00100000001000";
		Trees_din <= x"001f2035";
		wait for Clk_period;
		Addr <=  "00100000001001";
		Trees_din <= x"008e2035";
		wait for Clk_period;
		Addr <=  "00100000001010";
		Trees_din <= x"000e4f04";
		wait for Clk_period;
		Addr <=  "00100000001011";
		Trees_din <= x"005a2035";
		wait for Clk_period;
		Addr <=  "00100000001100";
		Trees_din <= x"ffa32035";
		wait for Clk_period;
		Addr <=  "00100000001101";
		Trees_din <= x"21000040";
		wait for Clk_period;
		Addr <=  "00100000001110";
		Trees_din <= x"21000038";
		wait for Clk_period;
		Addr <=  "00100000001111";
		Trees_din <= x"0109691c";
		wait for Clk_period;
		Addr <=  "00100000010000";
		Trees_din <= x"12037510";
		wait for Clk_period;
		Addr <=  "00100000010001";
		Trees_din <= x"12012308";
		wait for Clk_period;
		Addr <=  "00100000010010";
		Trees_din <= x"09005604";
		wait for Clk_period;
		Addr <=  "00100000010011";
		Trees_din <= x"ffc020e9";
		wait for Clk_period;
		Addr <=  "00100000010100";
		Trees_din <= x"001920e9";
		wait for Clk_period;
		Addr <=  "00100000010101";
		Trees_din <= x"05fde504";
		wait for Clk_period;
		Addr <=  "00100000010110";
		Trees_din <= x"002a20e9";
		wait for Clk_period;
		Addr <=  "00100000010111";
		Trees_din <= x"ff8820e9";
		wait for Clk_period;
		Addr <=  "00100000011000";
		Trees_din <= x"08030108";
		wait for Clk_period;
		Addr <=  "00100000011001";
		Trees_din <= x"1d005104";
		wait for Clk_period;
		Addr <=  "00100000011010";
		Trees_din <= x"ff7a20e9";
		wait for Clk_period;
		Addr <=  "00100000011011";
		Trees_din <= x"fffc20e9";
		wait for Clk_period;
		Addr <=  "00100000011100";
		Trees_din <= x"007020e9";
		wait for Clk_period;
		Addr <=  "00100000011101";
		Trees_din <= x"05fa3810";
		wait for Clk_period;
		Addr <=  "00100000011110";
		Trees_din <= x"020a7308";
		wait for Clk_period;
		Addr <=  "00100000011111";
		Trees_din <= x"0111ec04";
		wait for Clk_period;
		Addr <=  "00100000100000";
		Trees_din <= x"fff220e9";
		wait for Clk_period;
		Addr <=  "00100000100001";
		Trees_din <= x"003120e9";
		wait for Clk_period;
		Addr <=  "00100000100010";
		Trees_din <= x"0efd7604";
		wait for Clk_period;
		Addr <=  "00100000100011";
		Trees_din <= x"000f20e9";
		wait for Clk_period;
		Addr <=  "00100000100100";
		Trees_din <= x"ff8d20e9";
		wait for Clk_period;
		Addr <=  "00100000100101";
		Trees_din <= x"00153208";
		wait for Clk_period;
		Addr <=  "00100000100110";
		Trees_din <= x"04fb2804";
		wait for Clk_period;
		Addr <=  "00100000100111";
		Trees_din <= x"004b20e9";
		wait for Clk_period;
		Addr <=  "00100000101000";
		Trees_din <= x"000e20e9";
		wait for Clk_period;
		Addr <=  "00100000101001";
		Trees_din <= x"ff9620e9";
		wait for Clk_period;
		Addr <=  "00100000101010";
		Trees_din <= x"07005804";
		wait for Clk_period;
		Addr <=  "00100000101011";
		Trees_din <= x"001d20e9";
		wait for Clk_period;
		Addr <=  "00100000101100";
		Trees_din <= x"00bf20e9";
		wait for Clk_period;
		Addr <=  "00100000101101";
		Trees_din <= x"1403e418";
		wait for Clk_period;
		Addr <=  "00100000101110";
		Trees_din <= x"04fea40c";
		wait for Clk_period;
		Addr <=  "00100000101111";
		Trees_din <= x"03f2f604";
		wait for Clk_period;
		Addr <=  "00100000110000";
		Trees_din <= x"000920e9";
		wait for Clk_period;
		Addr <=  "00100000110001";
		Trees_din <= x"12026204";
		wait for Clk_period;
		Addr <=  "00100000110010";
		Trees_din <= x"ff6c20e9";
		wait for Clk_period;
		Addr <=  "00100000110011";
		Trees_din <= x"ffd820e9";
		wait for Clk_period;
		Addr <=  "00100000110100";
		Trees_din <= x"01074704";
		wait for Clk_period;
		Addr <=  "00100000110101";
		Trees_din <= x"ffac20e9";
		wait for Clk_period;
		Addr <=  "00100000110110";
		Trees_din <= x"0c015904";
		wait for Clk_period;
		Addr <=  "00100000110111";
		Trees_din <= x"006420e9";
		wait for Clk_period;
		Addr <=  "00100000111000";
		Trees_din <= x"ffed20e9";
		wait for Clk_period;
		Addr <=  "00100000111001";
		Trees_din <= x"006c20e9";
		wait for Clk_period;
		Addr <=  "00100000111010";
		Trees_din <= x"0c001910";
		wait for Clk_period;
		Addr <=  "00100000111011";
		Trees_din <= x"0e00880c";
		wait for Clk_period;
		Addr <=  "00100000111100";
		Trees_din <= x"06f9b608";
		wait for Clk_period;
		Addr <=  "00100000111101";
		Trees_din <= x"09005604";
		wait for Clk_period;
		Addr <=  "00100000111110";
		Trees_din <= x"00b22175";
		wait for Clk_period;
		Addr <=  "00100000111111";
		Trees_din <= x"00122175";
		wait for Clk_period;
		Addr <=  "00100001000000";
		Trees_din <= x"fffb2175";
		wait for Clk_period;
		Addr <=  "00100001000001";
		Trees_din <= x"ffb92175";
		wait for Clk_period;
		Addr <=  "00100001000010";
		Trees_din <= x"10f72510";
		wait for Clk_period;
		Addr <=  "00100001000011";
		Trees_din <= x"00042108";
		wait for Clk_period;
		Addr <=  "00100001000100";
		Trees_din <= x"0a02ad04";
		wait for Clk_period;
		Addr <=  "00100001000101";
		Trees_din <= x"001d2175";
		wait for Clk_period;
		Addr <=  "00100001000110";
		Trees_din <= x"00a02175";
		wait for Clk_period;
		Addr <=  "00100001000111";
		Trees_din <= x"010d9004";
		wait for Clk_period;
		Addr <=  "00100001001000";
		Trees_din <= x"ff8f2175";
		wait for Clk_period;
		Addr <=  "00100001001001";
		Trees_din <= x"005f2175";
		wait for Clk_period;
		Addr <=  "00100001001010";
		Trees_din <= x"1f001420";
		wait for Clk_period;
		Addr <=  "00100001001011";
		Trees_din <= x"01082a10";
		wait for Clk_period;
		Addr <=  "00100001001100";
		Trees_din <= x"07005d08";
		wait for Clk_period;
		Addr <=  "00100001001101";
		Trees_din <= x"0107ac04";
		wait for Clk_period;
		Addr <=  "00100001001110";
		Trees_din <= x"fff22175";
		wait for Clk_period;
		Addr <=  "00100001001111";
		Trees_din <= x"ff9a2175";
		wait for Clk_period;
		Addr <=  "00100001010000";
		Trees_din <= x"09005404";
		wait for Clk_period;
		Addr <=  "00100001010001";
		Trees_din <= x"00102175";
		wait for Clk_period;
		Addr <=  "00100001010010";
		Trees_din <= x"008b2175";
		wait for Clk_period;
		Addr <=  "00100001010011";
		Trees_din <= x"05fb9c08";
		wait for Clk_period;
		Addr <=  "00100001010100";
		Trees_din <= x"19008e04";
		wait for Clk_period;
		Addr <=  "00100001010101";
		Trees_din <= x"001c2175";
		wait for Clk_period;
		Addr <=  "00100001010110";
		Trees_din <= x"fff22175";
		wait for Clk_period;
		Addr <=  "00100001010111";
		Trees_din <= x"11012e04";
		wait for Clk_period;
		Addr <=  "00100001011000";
		Trees_din <= x"ffe12175";
		wait for Clk_period;
		Addr <=  "00100001011001";
		Trees_din <= x"00472175";
		wait for Clk_period;
		Addr <=  "00100001011010";
		Trees_din <= x"03fc9704";
		wait for Clk_period;
		Addr <=  "00100001011011";
		Trees_din <= x"ff7d2175";
		wait for Clk_period;
		Addr <=  "00100001011100";
		Trees_din <= x"001f2175";
		wait for Clk_period;
		Addr <=  "00100001011101";
		Trees_din <= x"0bf93224";
		wait for Clk_period;
		Addr <=  "00100001011110";
		Trees_din <= x"1c00371c";
		wait for Clk_period;
		Addr <=  "00100001011111";
		Trees_din <= x"1e006614";
		wait for Clk_period;
		Addr <=  "00100001100000";
		Trees_din <= x"1a00e108";
		wait for Clk_period;
		Addr <=  "00100001100001";
		Trees_din <= x"1b003304";
		wait for Clk_period;
		Addr <=  "00100001100010";
		Trees_din <= x"ffd62251";
		wait for Clk_period;
		Addr <=  "00100001100011";
		Trees_din <= x"ff792251";
		wait for Clk_period;
		Addr <=  "00100001100100";
		Trees_din <= x"01085b04";
		wait for Clk_period;
		Addr <=  "00100001100101";
		Trees_din <= x"ffa22251";
		wait for Clk_period;
		Addr <=  "00100001100110";
		Trees_din <= x"12011f04";
		wait for Clk_period;
		Addr <=  "00100001100111";
		Trees_din <= x"ffeb2251";
		wait for Clk_period;
		Addr <=  "00100001101000";
		Trees_din <= x"00882251";
		wait for Clk_period;
		Addr <=  "00100001101001";
		Trees_din <= x"06f4ba04";
		wait for Clk_period;
		Addr <=  "00100001101010";
		Trees_din <= x"00022251";
		wait for Clk_period;
		Addr <=  "00100001101011";
		Trees_din <= x"00aa2251";
		wait for Clk_period;
		Addr <=  "00100001101100";
		Trees_din <= x"02003504";
		wait for Clk_period;
		Addr <=  "00100001101101";
		Trees_din <= x"001a2251";
		wait for Clk_period;
		Addr <=  "00100001101110";
		Trees_din <= x"ff632251";
		wait for Clk_period;
		Addr <=  "00100001101111";
		Trees_din <= x"04f69f24";
		wait for Clk_period;
		Addr <=  "00100001110000";
		Trees_din <= x"1602d918";
		wait for Clk_period;
		Addr <=  "00100001110001";
		Trees_din <= x"1601030c";
		wait for Clk_period;
		Addr <=  "00100001110010";
		Trees_din <= x"0200af04";
		wait for Clk_period;
		Addr <=  "00100001110011";
		Trees_din <= x"00392251";
		wait for Clk_period;
		Addr <=  "00100001110100";
		Trees_din <= x"06fcc204";
		wait for Clk_period;
		Addr <=  "00100001110101";
		Trees_din <= x"ff7e2251";
		wait for Clk_period;
		Addr <=  "00100001110110";
		Trees_din <= x"ffdb2251";
		wait for Clk_period;
		Addr <=  "00100001110111";
		Trees_din <= x"1202ab08";
		wait for Clk_period;
		Addr <=  "00100001111000";
		Trees_din <= x"1500a004";
		wait for Clk_period;
		Addr <=  "00100001111001";
		Trees_din <= x"00732251";
		wait for Clk_period;
		Addr <=  "00100001111010";
		Trees_din <= x"ffd42251";
		wait for Clk_period;
		Addr <=  "00100001111011";
		Trees_din <= x"ffb52251";
		wait for Clk_period;
		Addr <=  "00100001111100";
		Trees_din <= x"09005a08";
		wait for Clk_period;
		Addr <=  "00100001111101";
		Trees_din <= x"05f70004";
		wait for Clk_period;
		Addr <=  "00100001111110";
		Trees_din <= x"00022251";
		wait for Clk_period;
		Addr <=  "00100001111111";
		Trees_din <= x"ff802251";
		wait for Clk_period;
		Addr <=  "00100010000000";
		Trees_din <= x"00202251";
		wait for Clk_period;
		Addr <=  "00100010000001";
		Trees_din <= x"03f31e0c";
		wait for Clk_period;
		Addr <=  "00100010000010";
		Trees_din <= x"06f30204";
		wait for Clk_period;
		Addr <=  "00100010000011";
		Trees_din <= x"ffc22251";
		wait for Clk_period;
		Addr <=  "00100010000100";
		Trees_din <= x"0c01ad04";
		wait for Clk_period;
		Addr <=  "00100010000101";
		Trees_din <= x"001c2251";
		wait for Clk_period;
		Addr <=  "00100010000110";
		Trees_din <= x"00c62251";
		wait for Clk_period;
		Addr <=  "00100010000111";
		Trees_din <= x"06fc3d10";
		wait for Clk_period;
		Addr <=  "00100010001000";
		Trees_din <= x"0d03ea08";
		wait for Clk_period;
		Addr <=  "00100010001001";
		Trees_din <= x"12028704";
		wait for Clk_period;
		Addr <=  "00100010001010";
		Trees_din <= x"000c2251";
		wait for Clk_period;
		Addr <=  "00100010001011";
		Trees_din <= x"ffed2251";
		wait for Clk_period;
		Addr <=  "00100010001100";
		Trees_din <= x"000b5604";
		wait for Clk_period;
		Addr <=  "00100010001101";
		Trees_din <= x"ffef2251";
		wait for Clk_period;
		Addr <=  "00100010001110";
		Trees_din <= x"ff7c2251";
		wait for Clk_period;
		Addr <=  "00100010001111";
		Trees_din <= x"01031d04";
		wait for Clk_period;
		Addr <=  "00100010010000";
		Trees_din <= x"ffef2251";
		wait for Clk_period;
		Addr <=  "00100010010001";
		Trees_din <= x"0f02dd04";
		wait for Clk_period;
		Addr <=  "00100010010010";
		Trees_din <= x"00702251";
		wait for Clk_period;
		Addr <=  "00100010010011";
		Trees_din <= x"ffed2251";
		wait for Clk_period;
		Addr <=  "00100010010100";
		Trees_din <= x"010d4f38";
		wait for Clk_period;
		Addr <=  "00100010010101";
		Trees_din <= x"03f6f418";
		wait for Clk_period;
		Addr <=  "00100010010110";
		Trees_din <= x"10028710";
		wait for Clk_period;
		Addr <=  "00100010010111";
		Trees_din <= x"14017204";
		wait for Clk_period;
		Addr <=  "00100010011000";
		Trees_din <= x"ffa8237d";
		wait for Clk_period;
		Addr <=  "00100010011001";
		Trees_din <= x"06f52304";
		wait for Clk_period;
		Addr <=  "00100010011010";
		Trees_din <= x"ffa9237d";
		wait for Clk_period;
		Addr <=  "00100010011011";
		Trees_din <= x"06f76d04";
		wait for Clk_period;
		Addr <=  "00100010011100";
		Trees_din <= x"0099237d";
		wait for Clk_period;
		Addr <=  "00100010011101";
		Trees_din <= x"ffd5237d";
		wait for Clk_period;
		Addr <=  "00100010011110";
		Trees_din <= x"04f58904";
		wait for Clk_period;
		Addr <=  "00100010011111";
		Trees_din <= x"ffda237d";
		wait for Clk_period;
		Addr <=  "00100010100000";
		Trees_din <= x"ff6d237d";
		wait for Clk_period;
		Addr <=  "00100010100001";
		Trees_din <= x"010d281c";
		wait for Clk_period;
		Addr <=  "00100010100010";
		Trees_din <= x"010cb410";
		wait for Clk_period;
		Addr <=  "00100010100011";
		Trees_din <= x"0c004108";
		wait for Clk_period;
		Addr <=  "00100010100100";
		Trees_din <= x"0d001a04";
		wait for Clk_period;
		Addr <=  "00100010100101";
		Trees_din <= x"ffe1237d";
		wait for Clk_period;
		Addr <=  "00100010100110";
		Trees_din <= x"005e237d";
		wait for Clk_period;
		Addr <=  "00100010100111";
		Trees_din <= x"0d00a704";
		wait for Clk_period;
		Addr <=  "00100010101000";
		Trees_din <= x"ffca237d";
		wait for Clk_period;
		Addr <=  "00100010101001";
		Trees_din <= x"0005237d";
		wait for Clk_period;
		Addr <=  "00100010101010";
		Trees_din <= x"18003704";
		wait for Clk_period;
		Addr <=  "00100010101011";
		Trees_din <= x"ff8d237d";
		wait for Clk_period;
		Addr <=  "00100010101100";
		Trees_din <= x"1c003804";
		wait for Clk_period;
		Addr <=  "00100010101101";
		Trees_din <= x"009f237d";
		wait for Clk_period;
		Addr <=  "00100010101110";
		Trees_din <= x"0013237d";
		wait for Clk_period;
		Addr <=  "00100010101111";
		Trees_din <= x"ff86237d";
		wait for Clk_period;
		Addr <=  "00100010110000";
		Trees_din <= x"0a028834";
		wait for Clk_period;
		Addr <=  "00100010110001";
		Trees_din <= x"1b00401c";
		wait for Clk_period;
		Addr <=  "00100010110010";
		Trees_din <= x"1e006a10";
		wait for Clk_period;
		Addr <=  "00100010110011";
		Trees_din <= x"000c5808";
		wait for Clk_period;
		Addr <=  "00100010110100";
		Trees_din <= x"09005904";
		wait for Clk_period;
		Addr <=  "00100010110101";
		Trees_din <= x"0061237d";
		wait for Clk_period;
		Addr <=  "00100010110110";
		Trees_din <= x"ffbc237d";
		wait for Clk_period;
		Addr <=  "00100010110111";
		Trees_din <= x"08030a04";
		wait for Clk_period;
		Addr <=  "00100010111000";
		Trees_din <= x"ffd5237d";
		wait for Clk_period;
		Addr <=  "00100010111001";
		Trees_din <= x"0073237d";
		wait for Clk_period;
		Addr <=  "00100010111010";
		Trees_din <= x"1d004204";
		wait for Clk_period;
		Addr <=  "00100010111011";
		Trees_din <= x"ff89237d";
		wait for Clk_period;
		Addr <=  "00100010111100";
		Trees_din <= x"1603f604";
		wait for Clk_period;
		Addr <=  "00100010111101";
		Trees_din <= x"0070237d";
		wait for Clk_period;
		Addr <=  "00100010111110";
		Trees_din <= x"ff9c237d";
		wait for Clk_period;
		Addr <=  "00100010111111";
		Trees_din <= x"06f5dc0c";
		wait for Clk_period;
		Addr <=  "00100011000000";
		Trees_din <= x"10fa3b04";
		wait for Clk_period;
		Addr <=  "00100011000001";
		Trees_din <= x"004b237d";
		wait for Clk_period;
		Addr <=  "00100011000010";
		Trees_din <= x"04ffda04";
		wait for Clk_period;
		Addr <=  "00100011000011";
		Trees_din <= x"ff89237d";
		wait for Clk_period;
		Addr <=  "00100011000100";
		Trees_din <= x"002c237d";
		wait for Clk_period;
		Addr <=  "00100011000101";
		Trees_din <= x"0800ea08";
		wait for Clk_period;
		Addr <=  "00100011000110";
		Trees_din <= x"08000d04";
		wait for Clk_period;
		Addr <=  "00100011000111";
		Trees_din <= x"ffe7237d";
		wait for Clk_period;
		Addr <=  "00100011001000";
		Trees_din <= x"0099237d";
		wait for Clk_period;
		Addr <=  "00100011001001";
		Trees_din <= x"ffaa237d";
		wait for Clk_period;
		Addr <=  "00100011001010";
		Trees_din <= x"1200de18";
		wait for Clk_period;
		Addr <=  "00100011001011";
		Trees_din <= x"0b03ba0c";
		wait for Clk_period;
		Addr <=  "00100011001100";
		Trees_din <= x"08030108";
		wait for Clk_period;
		Addr <=  "00100011001101";
		Trees_din <= x"18003f04";
		wait for Clk_period;
		Addr <=  "00100011001110";
		Trees_din <= x"001e237d";
		wait for Clk_period;
		Addr <=  "00100011001111";
		Trees_din <= x"0094237d";
		wait for Clk_period;
		Addr <=  "00100011010000";
		Trees_din <= x"ffc2237d";
		wait for Clk_period;
		Addr <=  "00100011010001";
		Trees_din <= x"000ae804";
		wait for Clk_period;
		Addr <=  "00100011010010";
		Trees_din <= x"0051237d";
		wait for Clk_period;
		Addr <=  "00100011010011";
		Trees_din <= x"0c02dd04";
		wait for Clk_period;
		Addr <=  "00100011010100";
		Trees_din <= x"ff8e237d";
		wait for Clk_period;
		Addr <=  "00100011010101";
		Trees_din <= x"0041237d";
		wait for Clk_period;
		Addr <=  "00100011010110";
		Trees_din <= x"1e008210";
		wait for Clk_period;
		Addr <=  "00100011010111";
		Trees_din <= x"17006c08";
		wait for Clk_period;
		Addr <=  "00100011011000";
		Trees_din <= x"1d003b04";
		wait for Clk_period;
		Addr <=  "00100011011001";
		Trees_din <= x"ffeb237d";
		wait for Clk_period;
		Addr <=  "00100011011010";
		Trees_din <= x"ff5d237d";
		wait for Clk_period;
		Addr <=  "00100011011011";
		Trees_din <= x"03f82f04";
		wait for Clk_period;
		Addr <=  "00100011011100";
		Trees_din <= x"ff9e237d";
		wait for Clk_period;
		Addr <=  "00100011011101";
		Trees_din <= x"0069237d";
		wait for Clk_period;
		Addr <=  "00100011011110";
		Trees_din <= x"006b237d";
		wait for Clk_period;
		Addr <=  "00100011011111";
		Trees_din <= x"1f000070";
		wait for Clk_period;
		Addr <=  "00100011100000";
		Trees_din <= x"010d4f30";
		wait for Clk_period;
		Addr <=  "00100011100001";
		Trees_din <= x"0010b11c";
		wait for Clk_period;
		Addr <=  "00100011100010";
		Trees_din <= x"0e02fe0c";
		wait for Clk_period;
		Addr <=  "00100011100011";
		Trees_din <= x"0e02d808";
		wait for Clk_period;
		Addr <=  "00100011100100";
		Trees_din <= x"15009904";
		wait for Clk_period;
		Addr <=  "00100011100101";
		Trees_din <= x"001c24b9";
		wait for Clk_period;
		Addr <=  "00100011100110";
		Trees_din <= x"ffec24b9";
		wait for Clk_period;
		Addr <=  "00100011100111";
		Trees_din <= x"00a924b9";
		wait for Clk_period;
		Addr <=  "00100011101000";
		Trees_din <= x"06f3d608";
		wait for Clk_period;
		Addr <=  "00100011101001";
		Trees_din <= x"1b003904";
		wait for Clk_period;
		Addr <=  "00100011101010";
		Trees_din <= x"007e24b9";
		wait for Clk_period;
		Addr <=  "00100011101011";
		Trees_din <= x"ffef24b9";
		wait for Clk_period;
		Addr <=  "00100011101100";
		Trees_din <= x"06f73004";
		wait for Clk_period;
		Addr <=  "00100011101101";
		Trees_din <= x"ff7c24b9";
		wait for Clk_period;
		Addr <=  "00100011101110";
		Trees_din <= x"ffec24b9";
		wait for Clk_period;
		Addr <=  "00100011101111";
		Trees_din <= x"1c003a10";
		wait for Clk_period;
		Addr <=  "00100011110000";
		Trees_din <= x"09005a08";
		wait for Clk_period;
		Addr <=  "00100011110001";
		Trees_din <= x"04fd5304";
		wait for Clk_period;
		Addr <=  "00100011110010";
		Trees_din <= x"ffbf24b9";
		wait for Clk_period;
		Addr <=  "00100011110011";
		Trees_din <= x"005d24b9";
		wait for Clk_period;
		Addr <=  "00100011110100";
		Trees_din <= x"1102fb04";
		wait for Clk_period;
		Addr <=  "00100011110101";
		Trees_din <= x"000324b9";
		wait for Clk_period;
		Addr <=  "00100011110110";
		Trees_din <= x"00c324b9";
		wait for Clk_period;
		Addr <=  "00100011110111";
		Trees_din <= x"ff7224b9";
		wait for Clk_period;
		Addr <=  "00100011111000";
		Trees_din <= x"13014820";
		wait for Clk_period;
		Addr <=  "00100011111001";
		Trees_din <= x"0a028810";
		wait for Clk_period;
		Addr <=  "00100011111010";
		Trees_din <= x"10056f08";
		wait for Clk_period;
		Addr <=  "00100011111011";
		Trees_din <= x"00119204";
		wait for Clk_period;
		Addr <=  "00100011111100";
		Trees_din <= x"003824b9";
		wait for Clk_period;
		Addr <=  "00100011111101";
		Trees_din <= x"ffef24b9";
		wait for Clk_period;
		Addr <=  "00100011111110";
		Trees_din <= x"03f97304";
		wait for Clk_period;
		Addr <=  "00100011111111";
		Trees_din <= x"ffb324b9";
		wait for Clk_period;
		Addr <=  "00100100000000";
		Trees_din <= x"004924b9";
		wait for Clk_period;
		Addr <=  "00100100000001";
		Trees_din <= x"18004c08";
		wait for Clk_period;
		Addr <=  "00100100000010";
		Trees_din <= x"17006c04";
		wait for Clk_period;
		Addr <=  "00100100000011";
		Trees_din <= x"ffa524b9";
		wait for Clk_period;
		Addr <=  "00100100000100";
		Trees_din <= x"001524b9";
		wait for Clk_period;
		Addr <=  "00100100000101";
		Trees_din <= x"0c016e04";
		wait for Clk_period;
		Addr <=  "00100100000110";
		Trees_din <= x"ffbf24b9";
		wait for Clk_period;
		Addr <=  "00100100000111";
		Trees_din <= x"008924b9";
		wait for Clk_period;
		Addr <=  "00100100001000";
		Trees_din <= x"010fff10";
		wait for Clk_period;
		Addr <=  "00100100001001";
		Trees_din <= x"06f83d08";
		wait for Clk_period;
		Addr <=  "00100100001010";
		Trees_din <= x"17012404";
		wait for Clk_period;
		Addr <=  "00100100001011";
		Trees_din <= x"00a224b9";
		wait for Clk_period;
		Addr <=  "00100100001100";
		Trees_din <= x"001b24b9";
		wait for Clk_period;
		Addr <=  "00100100001101";
		Trees_din <= x"08004904";
		wait for Clk_period;
		Addr <=  "00100100001110";
		Trees_din <= x"002b24b9";
		wait for Clk_period;
		Addr <=  "00100100001111";
		Trees_din <= x"ffb224b9";
		wait for Clk_period;
		Addr <=  "00100100010000";
		Trees_din <= x"0010d708";
		wait for Clk_period;
		Addr <=  "00100100010001";
		Trees_din <= x"0bfaee04";
		wait for Clk_period;
		Addr <=  "00100100010010";
		Trees_din <= x"ffcc24b9";
		wait for Clk_period;
		Addr <=  "00100100010011";
		Trees_din <= x"008b24b9";
		wait for Clk_period;
		Addr <=  "00100100010100";
		Trees_din <= x"0e03d004";
		wait for Clk_period;
		Addr <=  "00100100010101";
		Trees_din <= x"ff9b24b9";
		wait for Clk_period;
		Addr <=  "00100100010110";
		Trees_din <= x"000b24b9";
		wait for Clk_period;
		Addr <=  "00100100010111";
		Trees_din <= x"06f6f120";
		wait for Clk_period;
		Addr <=  "00100100011000";
		Trees_din <= x"0b04ee18";
		wait for Clk_period;
		Addr <=  "00100100011001";
		Trees_din <= x"0700580c";
		wait for Clk_period;
		Addr <=  "00100100011010";
		Trees_din <= x"1500af08";
		wait for Clk_period;
		Addr <=  "00100100011011";
		Trees_din <= x"0c037204";
		wait for Clk_period;
		Addr <=  "00100100011100";
		Trees_din <= x"ff6124b9";
		wait for Clk_period;
		Addr <=  "00100100011101";
		Trees_din <= x"001024b9";
		wait for Clk_period;
		Addr <=  "00100100011110";
		Trees_din <= x"002424b9";
		wait for Clk_period;
		Addr <=  "00100100011111";
		Trees_din <= x"1c003f08";
		wait for Clk_period;
		Addr <=  "00100100100000";
		Trees_din <= x"0afc8304";
		wait for Clk_period;
		Addr <=  "00100100100001";
		Trees_din <= x"003224b9";
		wait for Clk_period;
		Addr <=  "00100100100010";
		Trees_din <= x"ffb324b9";
		wait for Clk_period;
		Addr <=  "00100100100011";
		Trees_din <= x"006324b9";
		wait for Clk_period;
		Addr <=  "00100100100100";
		Trees_din <= x"18004004";
		wait for Clk_period;
		Addr <=  "00100100100101";
		Trees_din <= x"007824b9";
		wait for Clk_period;
		Addr <=  "00100100100110";
		Trees_din <= x"ffd924b9";
		wait for Clk_period;
		Addr <=  "00100100100111";
		Trees_din <= x"0f006a08";
		wait for Clk_period;
		Addr <=  "00100100101000";
		Trees_din <= x"00090504";
		wait for Clk_period;
		Addr <=  "00100100101001";
		Trees_din <= x"005e24b9";
		wait for Clk_period;
		Addr <=  "00100100101010";
		Trees_din <= x"ff8f24b9";
		wait for Clk_period;
		Addr <=  "00100100101011";
		Trees_din <= x"01082a04";
		wait for Clk_period;
		Addr <=  "00100100101100";
		Trees_din <= x"ffdb24b9";
		wait for Clk_period;
		Addr <=  "00100100101101";
		Trees_din <= x"00a024b9";
		wait for Clk_period;
		Addr <=  "00100100101110";
		Trees_din <= x"01fe6a04";
		wait for Clk_period;
		Addr <=  "00100100101111";
		Trees_din <= x"ff9e254d";
		wait for Clk_period;
		Addr <=  "00100100110000";
		Trees_din <= x"1500b22c";
		wait for Clk_period;
		Addr <=  "00100100110001";
		Trees_din <= x"1c002410";
		wait for Clk_period;
		Addr <=  "00100100110010";
		Trees_din <= x"02fffa04";
		wait for Clk_period;
		Addr <=  "00100100110011";
		Trees_din <= x"004e254d";
		wait for Clk_period;
		Addr <=  "00100100110100";
		Trees_din <= x"1401b104";
		wait for Clk_period;
		Addr <=  "00100100110101";
		Trees_din <= x"ff78254d";
		wait for Clk_period;
		Addr <=  "00100100110110";
		Trees_din <= x"0e01df04";
		wait for Clk_period;
		Addr <=  "00100100110111";
		Trees_din <= x"0005254d";
		wait for Clk_period;
		Addr <=  "00100100111000";
		Trees_din <= x"ffc5254d";
		wait for Clk_period;
		Addr <=  "00100100111001";
		Trees_din <= x"1703f610";
		wait for Clk_period;
		Addr <=  "00100100111010";
		Trees_din <= x"1603fa08";
		wait for Clk_period;
		Addr <=  "00100100111011";
		Trees_din <= x"07005e04";
		wait for Clk_period;
		Addr <=  "00100100111100";
		Trees_din <= x"0001254d";
		wait for Clk_period;
		Addr <=  "00100100111101";
		Trees_din <= x"0044254d";
		wait for Clk_period;
		Addr <=  "00100100111110";
		Trees_din <= x"1603ff04";
		wait for Clk_period;
		Addr <=  "00100100111111";
		Trees_din <= x"ffa5254d";
		wait for Clk_period;
		Addr <=  "00100101000000";
		Trees_din <= x"001e254d";
		wait for Clk_period;
		Addr <=  "00100101000001";
		Trees_din <= x"0d002a04";
		wait for Clk_period;
		Addr <=  "00100101000010";
		Trees_din <= x"ffd6254d";
		wait for Clk_period;
		Addr <=  "00100101000011";
		Trees_din <= x"04fc9804";
		wait for Clk_period;
		Addr <=  "00100101000100";
		Trees_din <= x"0019254d";
		wait for Clk_period;
		Addr <=  "00100101000101";
		Trees_din <= x"0088254d";
		wait for Clk_period;
		Addr <=  "00100101000110";
		Trees_din <= x"12027614";
		wait for Clk_period;
		Addr <=  "00100101000111";
		Trees_din <= x"0afb1808";
		wait for Clk_period;
		Addr <=  "00100101001000";
		Trees_din <= x"01094f04";
		wait for Clk_period;
		Addr <=  "00100101001001";
		Trees_din <= x"ffa7254d";
		wait for Clk_period;
		Addr <=  "00100101001010";
		Trees_din <= x"0028254d";
		wait for Clk_period;
		Addr <=  "00100101001011";
		Trees_din <= x"0e011708";
		wait for Clk_period;
		Addr <=  "00100101001100";
		Trees_din <= x"07005304";
		wait for Clk_period;
		Addr <=  "00100101001101";
		Trees_din <= x"ffab254d";
		wait for Clk_period;
		Addr <=  "00100101001110";
		Trees_din <= x"0062254d";
		wait for Clk_period;
		Addr <=  "00100101001111";
		Trees_din <= x"009f254d";
		wait for Clk_period;
		Addr <=  "00100101010000";
		Trees_din <= x"0c01bf04";
		wait for Clk_period;
		Addr <=  "00100101010001";
		Trees_din <= x"000b254d";
		wait for Clk_period;
		Addr <=  "00100101010010";
		Trees_din <= x"ff9b254d";
		wait for Clk_period;
		Addr <=  "00100101010011";
		Trees_din <= x"010f7450";
		wait for Clk_period;
		Addr <=  "00100101010100";
		Trees_din <= x"20040020";
		wait for Clk_period;
		Addr <=  "00100101010101";
		Trees_din <= x"09005a14";
		wait for Clk_period;
		Addr <=  "00100101010110";
		Trees_din <= x"05f86604";
		wait for Clk_period;
		Addr <=  "00100101010111";
		Trees_din <= x"00272659";
		wait for Clk_period;
		Addr <=  "00100101011000";
		Trees_din <= x"19008008";
		wait for Clk_period;
		Addr <=  "00100101011001";
		Trees_din <= x"18005104";
		wait for Clk_period;
		Addr <=  "00100101011010";
		Trees_din <= x"004e2659";
		wait for Clk_period;
		Addr <=  "00100101011011";
		Trees_din <= x"ffb82659";
		wait for Clk_period;
		Addr <=  "00100101011100";
		Trees_din <= x"1103fb04";
		wait for Clk_period;
		Addr <=  "00100101011101";
		Trees_din <= x"ff742659";
		wait for Clk_period;
		Addr <=  "00100101011110";
		Trees_din <= x"00172659";
		wait for Clk_period;
		Addr <=  "00100101011111";
		Trees_din <= x"10028708";
		wait for Clk_period;
		Addr <=  "00100101100000";
		Trees_din <= x"06f69e04";
		wait for Clk_period;
		Addr <=  "00100101100001";
		Trees_din <= x"00182659";
		wait for Clk_period;
		Addr <=  "00100101100010";
		Trees_din <= x"ff9d2659";
		wait for Clk_period;
		Addr <=  "00100101100011";
		Trees_din <= x"00862659";
		wait for Clk_period;
		Addr <=  "00100101100100";
		Trees_din <= x"1400b114";
		wait for Clk_period;
		Addr <=  "00100101100101";
		Trees_din <= x"1400a50c";
		wait for Clk_period;
		Addr <=  "00100101100110";
		Trees_din <= x"0e03ed08";
		wait for Clk_period;
		Addr <=  "00100101100111";
		Trees_din <= x"05f9de04";
		wait for Clk_period;
		Addr <=  "00100101101000";
		Trees_din <= x"ffbb2659";
		wait for Clk_period;
		Addr <=  "00100101101001";
		Trees_din <= x"00102659";
		wait for Clk_period;
		Addr <=  "00100101101010";
		Trees_din <= x"ff792659";
		wait for Clk_period;
		Addr <=  "00100101101011";
		Trees_din <= x"04004504";
		wait for Clk_period;
		Addr <=  "00100101101100";
		Trees_din <= x"ff712659";
		wait for Clk_period;
		Addr <=  "00100101101101";
		Trees_din <= x"ffde2659";
		wait for Clk_period;
		Addr <=  "00100101101110";
		Trees_din <= x"1400eb0c";
		wait for Clk_period;
		Addr <=  "00100101101111";
		Trees_din <= x"0f000304";
		wait for Clk_period;
		Addr <=  "00100101110000";
		Trees_din <= x"00a82659";
		wait for Clk_period;
		Addr <=  "00100101110001";
		Trees_din <= x"06f64804";
		wait for Clk_period;
		Addr <=  "00100101110010";
		Trees_din <= x"ffe02659";
		wait for Clk_period;
		Addr <=  "00100101110011";
		Trees_din <= x"00482659";
		wait for Clk_period;
		Addr <=  "00100101110100";
		Trees_din <= x"0f000f08";
		wait for Clk_period;
		Addr <=  "00100101110101";
		Trees_din <= x"04f81504";
		wait for Clk_period;
		Addr <=  "00100101110110";
		Trees_din <= x"00552659";
		wait for Clk_period;
		Addr <=  "00100101110111";
		Trees_din <= x"ff952659";
		wait for Clk_period;
		Addr <=  "00100101111000";
		Trees_din <= x"14010804";
		wait for Clk_period;
		Addr <=  "00100101111001";
		Trees_din <= x"ffab2659";
		wait for Clk_period;
		Addr <=  "00100101111010";
		Trees_din <= x"000c2659";
		wait for Clk_period;
		Addr <=  "00100101111011";
		Trees_din <= x"03f9f228";
		wait for Clk_period;
		Addr <=  "00100101111100";
		Trees_din <= x"21000020";
		wait for Clk_period;
		Addr <=  "00100101111101";
		Trees_din <= x"0b049d10";
		wait for Clk_period;
		Addr <=  "00100101111110";
		Trees_din <= x"0c00aa08";
		wait for Clk_period;
		Addr <=  "00100101111111";
		Trees_din <= x"1101fb04";
		wait for Clk_period;
		Addr <=  "00100110000000";
		Trees_din <= x"ffeb2659";
		wait for Clk_period;
		Addr <=  "00100110000001";
		Trees_din <= x"007d2659";
		wait for Clk_period;
		Addr <=  "00100110000010";
		Trees_din <= x"17001a04";
		wait for Clk_period;
		Addr <=  "00100110000011";
		Trees_din <= x"00162659";
		wait for Clk_period;
		Addr <=  "00100110000100";
		Trees_din <= x"ffc62659";
		wait for Clk_period;
		Addr <=  "00100110000101";
		Trees_din <= x"12febb08";
		wait for Clk_period;
		Addr <=  "00100110000110";
		Trees_din <= x"03f5dd04";
		wait for Clk_period;
		Addr <=  "00100110000111";
		Trees_din <= x"ff9f2659";
		wait for Clk_period;
		Addr <=  "00100110001000";
		Trees_din <= x"003e2659";
		wait for Clk_period;
		Addr <=  "00100110001001";
		Trees_din <= x"05fa0504";
		wait for Clk_period;
		Addr <=  "00100110001010";
		Trees_din <= x"008f2659";
		wait for Clk_period;
		Addr <=  "00100110001011";
		Trees_din <= x"00192659";
		wait for Clk_period;
		Addr <=  "00100110001100";
		Trees_din <= x"01128f04";
		wait for Clk_period;
		Addr <=  "00100110001101";
		Trees_din <= x"ff652659";
		wait for Clk_period;
		Addr <=  "00100110001110";
		Trees_din <= x"00072659";
		wait for Clk_period;
		Addr <=  "00100110001111";
		Trees_din <= x"0efa1a04";
		wait for Clk_period;
		Addr <=  "00100110010000";
		Trees_din <= x"ffee2659";
		wait for Clk_period;
		Addr <=  "00100110010001";
		Trees_din <= x"08001404";
		wait for Clk_period;
		Addr <=  "00100110010010";
		Trees_din <= x"fffe2659";
		wait for Clk_period;
		Addr <=  "00100110010011";
		Trees_din <= x"0d038804";
		wait for Clk_period;
		Addr <=  "00100110010100";
		Trees_din <= x"008d2659";
		wait for Clk_period;
		Addr <=  "00100110010101";
		Trees_din <= x"00202659";
		wait for Clk_period;
		Addr <=  "00100110010110";
		Trees_din <= x"1c004550";
		wait for Clk_period;
		Addr <=  "00100110010111";
		Trees_din <= x"18004818";
		wait for Clk_period;
		Addr <=  "00100110011000";
		Trees_din <= x"1d004d10";
		wait for Clk_period;
		Addr <=  "00100110011001";
		Trees_din <= x"1d004c0c";
		wait for Clk_period;
		Addr <=  "00100110011010";
		Trees_din <= x"1d004c08";
		wait for Clk_period;
		Addr <=  "00100110011011";
		Trees_din <= x"14027504";
		wait for Clk_period;
		Addr <=  "00100110011100";
		Trees_din <= x"0009275d";
		wait for Clk_period;
		Addr <=  "00100110011101";
		Trees_din <= x"ffea275d";
		wait for Clk_period;
		Addr <=  "00100110011110";
		Trees_din <= x"ff7b275d";
		wait for Clk_period;
		Addr <=  "00100110011111";
		Trees_din <= x"0089275d";
		wait for Clk_period;
		Addr <=  "00100110100000";
		Trees_din <= x"0f038a04";
		wait for Clk_period;
		Addr <=  "00100110100001";
		Trees_din <= x"ff7e275d";
		wait for Clk_period;
		Addr <=  "00100110100010";
		Trees_din <= x"000e275d";
		wait for Clk_period;
		Addr <=  "00100110100011";
		Trees_din <= x"02021b18";
		wait for Clk_period;
		Addr <=  "00100110100100";
		Trees_din <= x"010a420c";
		wait for Clk_period;
		Addr <=  "00100110100101";
		Trees_din <= x"0afb0104";
		wait for Clk_period;
		Addr <=  "00100110100110";
		Trees_din <= x"ffa5275d";
		wait for Clk_period;
		Addr <=  "00100110100111";
		Trees_din <= x"1a00b304";
		wait for Clk_period;
		Addr <=  "00100110101000";
		Trees_din <= x"0058275d";
		wait for Clk_period;
		Addr <=  "00100110101001";
		Trees_din <= x"ffd8275d";
		wait for Clk_period;
		Addr <=  "00100110101010";
		Trees_din <= x"00126b04";
		wait for Clk_period;
		Addr <=  "00100110101011";
		Trees_din <= x"0093275d";
		wait for Clk_period;
		Addr <=  "00100110101100";
		Trees_din <= x"13001304";
		wait for Clk_period;
		Addr <=  "00100110101101";
		Trees_din <= x"ffcf275d";
		wait for Clk_period;
		Addr <=  "00100110101110";
		Trees_din <= x"006f275d";
		wait for Clk_period;
		Addr <=  "00100110101111";
		Trees_din <= x"1a00ac10";
		wait for Clk_period;
		Addr <=  "00100110110000";
		Trees_din <= x"18004d08";
		wait for Clk_period;
		Addr <=  "00100110110001";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00100110110010";
		Trees_din <= x"fff0275d";
		wait for Clk_period;
		Addr <=  "00100110110011";
		Trees_din <= x"ff85275d";
		wait for Clk_period;
		Addr <=  "00100110110100";
		Trees_din <= x"04fdef04";
		wait for Clk_period;
		Addr <=  "00100110110101";
		Trees_din <= x"0050275d";
		wait for Clk_period;
		Addr <=  "00100110110110";
		Trees_din <= x"ffb3275d";
		wait for Clk_period;
		Addr <=  "00100110110111";
		Trees_din <= x"01096908";
		wait for Clk_period;
		Addr <=  "00100110111000";
		Trees_din <= x"1004d504";
		wait for Clk_period;
		Addr <=  "00100110111001";
		Trees_din <= x"ff8a275d";
		wait for Clk_period;
		Addr <=  "00100110111010";
		Trees_din <= x"0045275d";
		wait for Clk_period;
		Addr <=  "00100110111011";
		Trees_din <= x"10f97c04";
		wait for Clk_period;
		Addr <=  "00100110111100";
		Trees_din <= x"ffce275d";
		wait for Clk_period;
		Addr <=  "00100110111101";
		Trees_din <= x"006e275d";
		wait for Clk_period;
		Addr <=  "00100110111110";
		Trees_din <= x"04f8ba10";
		wait for Clk_period;
		Addr <=  "00100110111111";
		Trees_din <= x"13ff4408";
		wait for Clk_period;
		Addr <=  "00100111000000";
		Trees_din <= x"0c01e704";
		wait for Clk_period;
		Addr <=  "00100111000001";
		Trees_din <= x"ffe6275d";
		wait for Clk_period;
		Addr <=  "00100111000010";
		Trees_din <= x"0091275d";
		wait for Clk_period;
		Addr <=  "00100111000011";
		Trees_din <= x"16026704";
		wait for Clk_period;
		Addr <=  "00100111000100";
		Trees_din <= x"ffa9275d";
		wait for Clk_period;
		Addr <=  "00100111000101";
		Trees_din <= x"fffd275d";
		wait for Clk_period;
		Addr <=  "00100111000110";
		Trees_din <= x"0010d720";
		wait for Clk_period;
		Addr <=  "00100111000111";
		Trees_din <= x"03fae610";
		wait for Clk_period;
		Addr <=  "00100111001000";
		Trees_din <= x"06f5b408";
		wait for Clk_period;
		Addr <=  "00100111001001";
		Trees_din <= x"1a009a04";
		wait for Clk_period;
		Addr <=  "00100111001010";
		Trees_din <= x"007b275d";
		wait for Clk_period;
		Addr <=  "00100111001011";
		Trees_din <= x"ffd6275d";
		wait for Clk_period;
		Addr <=  "00100111001100";
		Trees_din <= x"010c6804";
		wait for Clk_period;
		Addr <=  "00100111001101";
		Trees_din <= x"ff8d275d";
		wait for Clk_period;
		Addr <=  "00100111001110";
		Trees_din <= x"000c275d";
		wait for Clk_period;
		Addr <=  "00100111001111";
		Trees_din <= x"03fee208";
		wait for Clk_period;
		Addr <=  "00100111010000";
		Trees_din <= x"1c004b04";
		wait for Clk_period;
		Addr <=  "00100111010001";
		Trees_din <= x"ff54275d";
		wait for Clk_period;
		Addr <=  "00100111010010";
		Trees_din <= x"fff6275d";
		wait for Clk_period;
		Addr <=  "00100111010011";
		Trees_din <= x"0afce404";
		wait for Clk_period;
		Addr <=  "00100111010100";
		Trees_din <= x"ffa8275d";
		wait for Clk_period;
		Addr <=  "00100111010101";
		Trees_din <= x"0040275d";
		wait for Clk_period;
		Addr <=  "00100111010110";
		Trees_din <= x"ff77275d";
		wait for Clk_period;
		Addr <=  "00100111010111";
		Trees_din <= x"0118036c";
		wait for Clk_period;
		Addr <=  "00100111011000";
		Trees_din <= x"15008330";
		wait for Clk_period;
		Addr <=  "00100111011001";
		Trees_din <= x"18004f14";
		wait for Clk_period;
		Addr <=  "00100111011010";
		Trees_din <= x"1402d208";
		wait for Clk_period;
		Addr <=  "00100111011011";
		Trees_din <= x"06f35804";
		wait for Clk_period;
		Addr <=  "00100111011100";
		Trees_din <= x"fff12839";
		wait for Clk_period;
		Addr <=  "00100111011101";
		Trees_din <= x"ff6b2839";
		wait for Clk_period;
		Addr <=  "00100111011110";
		Trees_din <= x"07004c04";
		wait for Clk_period;
		Addr <=  "00100111011111";
		Trees_din <= x"006f2839";
		wait for Clk_period;
		Addr <=  "00100111100000";
		Trees_din <= x"010d9004";
		wait for Clk_period;
		Addr <=  "00100111100001";
		Trees_din <= x"ff982839";
		wait for Clk_period;
		Addr <=  "00100111100010";
		Trees_din <= x"00292839";
		wait for Clk_period;
		Addr <=  "00100111100011";
		Trees_din <= x"0b03e310";
		wait for Clk_period;
		Addr <=  "00100111100100";
		Trees_din <= x"03fae608";
		wait for Clk_period;
		Addr <=  "00100111100101";
		Trees_din <= x"15007804";
		wait for Clk_period;
		Addr <=  "00100111100110";
		Trees_din <= x"ffd02839";
		wait for Clk_period;
		Addr <=  "00100111100111";
		Trees_din <= x"004f2839";
		wait for Clk_period;
		Addr <=  "00100111101000";
		Trees_din <= x"0f03ea04";
		wait for Clk_period;
		Addr <=  "00100111101001";
		Trees_din <= x"ff802839";
		wait for Clk_period;
		Addr <=  "00100111101010";
		Trees_din <= x"000f2839";
		wait for Clk_period;
		Addr <=  "00100111101011";
		Trees_din <= x"08000904";
		wait for Clk_period;
		Addr <=  "00100111101100";
		Trees_din <= x"ffb72839";
		wait for Clk_period;
		Addr <=  "00100111101101";
		Trees_din <= x"03f85a04";
		wait for Clk_period;
		Addr <=  "00100111101110";
		Trees_din <= x"fff42839";
		wait for Clk_period;
		Addr <=  "00100111101111";
		Trees_din <= x"00852839";
		wait for Clk_period;
		Addr <=  "00100111110000";
		Trees_din <= x"18004820";
		wait for Clk_period;
		Addr <=  "00100111110001";
		Trees_din <= x"0af7ba10";
		wait for Clk_period;
		Addr <=  "00100111110010";
		Trees_din <= x"19009108";
		wait for Clk_period;
		Addr <=  "00100111110011";
		Trees_din <= x"1603dd04";
		wait for Clk_period;
		Addr <=  "00100111110100";
		Trees_din <= x"009a2839";
		wait for Clk_period;
		Addr <=  "00100111110101";
		Trees_din <= x"00252839";
		wait for Clk_period;
		Addr <=  "00100111110110";
		Trees_din <= x"01094f04";
		wait for Clk_period;
		Addr <=  "00100111110111";
		Trees_din <= x"ffad2839";
		wait for Clk_period;
		Addr <=  "00100111111000";
		Trees_din <= x"003c2839";
		wait for Clk_period;
		Addr <=  "00100111111001";
		Trees_din <= x"0af7f108";
		wait for Clk_period;
		Addr <=  "00100111111010";
		Trees_din <= x"1703d804";
		wait for Clk_period;
		Addr <=  "00100111111011";
		Trees_din <= x"ff8d2839";
		wait for Clk_period;
		Addr <=  "00100111111100";
		Trees_din <= x"00302839";
		wait for Clk_period;
		Addr <=  "00100111111101";
		Trees_din <= x"15008f04";
		wait for Clk_period;
		Addr <=  "00100111111110";
		Trees_din <= x"ffd12839";
		wait for Clk_period;
		Addr <=  "00100111111111";
		Trees_din <= x"00022839";
		wait for Clk_period;
		Addr <=  "00101000000000";
		Trees_din <= x"02021b0c";
		wait for Clk_period;
		Addr <=  "00101000000001";
		Trees_din <= x"08016008";
		wait for Clk_period;
		Addr <=  "00101000000010";
		Trees_din <= x"06f38c04";
		wait for Clk_period;
		Addr <=  "00101000000011";
		Trees_din <= x"ffda2839";
		wait for Clk_period;
		Addr <=  "00101000000100";
		Trees_din <= x"00652839";
		wait for Clk_period;
		Addr <=  "00101000000101";
		Trees_din <= x"ffde2839";
		wait for Clk_period;
		Addr <=  "00101000000110";
		Trees_din <= x"1a00ac08";
		wait for Clk_period;
		Addr <=  "00101000000111";
		Trees_din <= x"1e008104";
		wait for Clk_period;
		Addr <=  "00101000001000";
		Trees_din <= x"ff9d2839";
		wait for Clk_period;
		Addr <=  "00101000001001";
		Trees_din <= x"00202839";
		wait for Clk_period;
		Addr <=  "00101000001010";
		Trees_din <= x"01090e04";
		wait for Clk_period;
		Addr <=  "00101000001011";
		Trees_din <= x"ffc92839";
		wait for Clk_period;
		Addr <=  "00101000001100";
		Trees_din <= x"00572839";
		wait for Clk_period;
		Addr <=  "00101000001101";
		Trees_din <= x"005d2839";
		wait for Clk_period;
		Addr <=  "00101000001110";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00101000001111";
		Trees_din <= x"01082a44";
		wait for Clk_period;
		Addr <=  "00101000010000";
		Trees_din <= x"07005d3c";
		wait for Clk_period;
		Addr <=  "00101000010001";
		Trees_din <= x"1200f71c";
		wait for Clk_period;
		Addr <=  "00101000010010";
		Trees_din <= x"05fe9610";
		wait for Clk_period;
		Addr <=  "00101000010011";
		Trees_din <= x"04f92008";
		wait for Clk_period;
		Addr <=  "00101000010100";
		Trees_din <= x"13fd6f04";
		wait for Clk_period;
		Addr <=  "00101000010101";
		Trees_din <= x"00412959";
		wait for Clk_period;
		Addr <=  "00101000010110";
		Trees_din <= x"ffb82959";
		wait for Clk_period;
		Addr <=  "00101000010111";
		Trees_din <= x"07004a04";
		wait for Clk_period;
		Addr <=  "00101000011000";
		Trees_din <= x"00392959";
		wait for Clk_period;
		Addr <=  "00101000011001";
		Trees_din <= x"ff952959";
		wait for Clk_period;
		Addr <=  "00101000011010";
		Trees_din <= x"0a019904";
		wait for Clk_period;
		Addr <=  "00101000011011";
		Trees_din <= x"ffd02959";
		wait for Clk_period;
		Addr <=  "00101000011100";
		Trees_din <= x"1a00ba04";
		wait for Clk_period;
		Addr <=  "00101000011101";
		Trees_din <= x"ffed2959";
		wait for Clk_period;
		Addr <=  "00101000011110";
		Trees_din <= x"007c2959";
		wait for Clk_period;
		Addr <=  "00101000011111";
		Trees_din <= x"1c003c10";
		wait for Clk_period;
		Addr <=  "00101000100000";
		Trees_din <= x"1d004408";
		wait for Clk_period;
		Addr <=  "00101000100001";
		Trees_din <= x"06f40d04";
		wait for Clk_period;
		Addr <=  "00101000100010";
		Trees_din <= x"00452959";
		wait for Clk_period;
		Addr <=  "00101000100011";
		Trees_din <= x"ffd62959";
		wait for Clk_period;
		Addr <=  "00101000100100";
		Trees_din <= x"13014104";
		wait for Clk_period;
		Addr <=  "00101000100101";
		Trees_din <= x"00742959";
		wait for Clk_period;
		Addr <=  "00101000100110";
		Trees_din <= x"ffad2959";
		wait for Clk_period;
		Addr <=  "00101000100111";
		Trees_din <= x"0f002c08";
		wait for Clk_period;
		Addr <=  "00101000101000";
		Trees_din <= x"05fb4504";
		wait for Clk_period;
		Addr <=  "00101000101001";
		Trees_din <= x"00572959";
		wait for Clk_period;
		Addr <=  "00101000101010";
		Trees_din <= x"ffe52959";
		wait for Clk_period;
		Addr <=  "00101000101011";
		Trees_din <= x"03029104";
		wait for Clk_period;
		Addr <=  "00101000101100";
		Trees_din <= x"ff742959";
		wait for Clk_period;
		Addr <=  "00101000101101";
		Trees_din <= x"fff32959";
		wait for Clk_period;
		Addr <=  "00101000101110";
		Trees_din <= x"19008804";
		wait for Clk_period;
		Addr <=  "00101000101111";
		Trees_din <= x"00722959";
		wait for Clk_period;
		Addr <=  "00101000110000";
		Trees_din <= x"00082959";
		wait for Clk_period;
		Addr <=  "00101000110001";
		Trees_din <= x"1900b034";
		wait for Clk_period;
		Addr <=  "00101000110010";
		Trees_din <= x"0bf95614";
		wait for Clk_period;
		Addr <=  "00101000110011";
		Trees_din <= x"0900570c";
		wait for Clk_period;
		Addr <=  "00101000110100";
		Trees_din <= x"1603e308";
		wait for Clk_period;
		Addr <=  "00101000110101";
		Trees_din <= x"10055404";
		wait for Clk_period;
		Addr <=  "00101000110110";
		Trees_din <= x"00372959";
		wait for Clk_period;
		Addr <=  "00101000110111";
		Trees_din <= x"ffab2959";
		wait for Clk_period;
		Addr <=  "00101000111000";
		Trees_din <= x"ffa12959";
		wait for Clk_period;
		Addr <=  "00101000111001";
		Trees_din <= x"17000204";
		wait for Clk_period;
		Addr <=  "00101000111010";
		Trees_din <= x"fff82959";
		wait for Clk_period;
		Addr <=  "00101000111011";
		Trees_din <= x"ff772959";
		wait for Clk_period;
		Addr <=  "00101000111100";
		Trees_din <= x"0bf99810";
		wait for Clk_period;
		Addr <=  "00101000111101";
		Trees_din <= x"1c003308";
		wait for Clk_period;
		Addr <=  "00101000111110";
		Trees_din <= x"07005604";
		wait for Clk_period;
		Addr <=  "00101000111111";
		Trees_din <= x"ffa72959";
		wait for Clk_period;
		Addr <=  "00101001000000";
		Trees_din <= x"00182959";
		wait for Clk_period;
		Addr <=  "00101001000001";
		Trees_din <= x"04041b04";
		wait for Clk_period;
		Addr <=  "00101001000010";
		Trees_din <= x"00832959";
		wait for Clk_period;
		Addr <=  "00101001000011";
		Trees_din <= x"ffd72959";
		wait for Clk_period;
		Addr <=  "00101001000100";
		Trees_din <= x"0f02d608";
		wait for Clk_period;
		Addr <=  "00101001000101";
		Trees_din <= x"1c002c04";
		wait for Clk_period;
		Addr <=  "00101001000110";
		Trees_din <= x"ffe22959";
		wait for Clk_period;
		Addr <=  "00101001000111";
		Trees_din <= x"00162959";
		wait for Clk_period;
		Addr <=  "00101001001000";
		Trees_din <= x"0c026304";
		wait for Clk_period;
		Addr <=  "00101001001001";
		Trees_din <= x"fff62959";
		wait for Clk_period;
		Addr <=  "00101001001010";
		Trees_din <= x"ff862959";
		wait for Clk_period;
		Addr <=  "00101001001011";
		Trees_din <= x"11009008";
		wait for Clk_period;
		Addr <=  "00101001001100";
		Trees_din <= x"02062104";
		wait for Clk_period;
		Addr <=  "00101001001101";
		Trees_din <= x"000d2959";
		wait for Clk_period;
		Addr <=  "00101001001110";
		Trees_din <= x"ff992959";
		wait for Clk_period;
		Addr <=  "00101001001111";
		Trees_din <= x"0011570c";
		wait for Clk_period;
		Addr <=  "00101001010000";
		Trees_din <= x"07004f04";
		wait for Clk_period;
		Addr <=  "00101001010001";
		Trees_din <= x"00082959";
		wait for Clk_period;
		Addr <=  "00101001010010";
		Trees_din <= x"14026e04";
		wait for Clk_period;
		Addr <=  "00101001010011";
		Trees_din <= x"00a22959";
		wait for Clk_period;
		Addr <=  "00101001010100";
		Trees_din <= x"002a2959";
		wait for Clk_period;
		Addr <=  "00101001010101";
		Trees_din <= x"ffc02959";
		wait for Clk_period;
		Addr <=  "00101001010110";
		Trees_din <= x"010cb468";
		wait for Clk_period;
		Addr <=  "00101001010111";
		Trees_din <= x"1400b128";
		wait for Clk_period;
		Addr <=  "00101001011000";
		Trees_din <= x"1400871c";
		wait for Clk_period;
		Addr <=  "00101001011001";
		Trees_din <= x"0e01d610";
		wait for Clk_period;
		Addr <=  "00101001011010";
		Trees_din <= x"1003dd08";
		wait for Clk_period;
		Addr <=  "00101001011011";
		Trees_din <= x"0b03ba04";
		wait for Clk_period;
		Addr <=  "00101001011100";
		Trees_din <= x"00082ad5";
		wait for Clk_period;
		Addr <=  "00101001011101";
		Trees_din <= x"ff802ad5";
		wait for Clk_period;
		Addr <=  "00101001011110";
		Trees_din <= x"12fe4404";
		wait for Clk_period;
		Addr <=  "00101001011111";
		Trees_din <= x"ffaf2ad5";
		wait for Clk_period;
		Addr <=  "00101001100000";
		Trees_din <= x"00402ad5";
		wait for Clk_period;
		Addr <=  "00101001100001";
		Trees_din <= x"07005204";
		wait for Clk_period;
		Addr <=  "00101001100010";
		Trees_din <= x"000f2ad5";
		wait for Clk_period;
		Addr <=  "00101001100011";
		Trees_din <= x"10f9ef04";
		wait for Clk_period;
		Addr <=  "00101001100100";
		Trees_din <= x"000c2ad5";
		wait for Clk_period;
		Addr <=  "00101001100101";
		Trees_din <= x"ff792ad5";
		wait for Clk_period;
		Addr <=  "00101001100110";
		Trees_din <= x"1500a204";
		wait for Clk_period;
		Addr <=  "00101001100111";
		Trees_din <= x"ff702ad5";
		wait for Clk_period;
		Addr <=  "00101001101000";
		Trees_din <= x"04fe1204";
		wait for Clk_period;
		Addr <=  "00101001101001";
		Trees_din <= x"ff8f2ad5";
		wait for Clk_period;
		Addr <=  "00101001101010";
		Trees_din <= x"00452ad5";
		wait for Clk_period;
		Addr <=  "00101001101011";
		Trees_din <= x"14028020";
		wait for Clk_period;
		Addr <=  "00101001101100";
		Trees_din <= x"07005a10";
		wait for Clk_period;
		Addr <=  "00101001101101";
		Trees_din <= x"01084108";
		wait for Clk_period;
		Addr <=  "00101001101110";
		Trees_din <= x"03faba04";
		wait for Clk_period;
		Addr <=  "00101001101111";
		Trees_din <= x"ffae2ad5";
		wait for Clk_period;
		Addr <=  "00101001110000";
		Trees_din <= x"00112ad5";
		wait for Clk_period;
		Addr <=  "00101001110001";
		Trees_din <= x"1500a004";
		wait for Clk_period;
		Addr <=  "00101001110010";
		Trees_din <= x"005b2ad5";
		wait for Clk_period;
		Addr <=  "00101001110011";
		Trees_din <= x"ffe82ad5";
		wait for Clk_period;
		Addr <=  "00101001110100";
		Trees_din <= x"1003dd08";
		wait for Clk_period;
		Addr <=  "00101001110101";
		Trees_din <= x"0e03b204";
		wait for Clk_period;
		Addr <=  "00101001110110";
		Trees_din <= x"ff822ad5";
		wait for Clk_period;
		Addr <=  "00101001110111";
		Trees_din <= x"001c2ad5";
		wait for Clk_period;
		Addr <=  "00101001111000";
		Trees_din <= x"0003aa04";
		wait for Clk_period;
		Addr <=  "00101001111001";
		Trees_din <= x"ffa22ad5";
		wait for Clk_period;
		Addr <=  "00101001111010";
		Trees_din <= x"00442ad5";
		wait for Clk_period;
		Addr <=  "00101001111011";
		Trees_din <= x"14032e10";
		wait for Clk_period;
		Addr <=  "00101001111100";
		Trees_din <= x"1b003708";
		wait for Clk_period;
		Addr <=  "00101001111101";
		Trees_din <= x"1b003504";
		wait for Clk_period;
		Addr <=  "00101001111110";
		Trees_din <= x"ffd22ad5";
		wait for Clk_period;
		Addr <=  "00101001111111";
		Trees_din <= x"00792ad5";
		wait for Clk_period;
		Addr <=  "00101010000000";
		Trees_din <= x"00011804";
		wait for Clk_period;
		Addr <=  "00101010000001";
		Trees_din <= x"ffd92ad5";
		wait for Clk_period;
		Addr <=  "00101010000010";
		Trees_din <= x"ff612ad5";
		wait for Clk_period;
		Addr <=  "00101010000011";
		Trees_din <= x"09005808";
		wait for Clk_period;
		Addr <=  "00101010000100";
		Trees_din <= x"0c01c804";
		wait for Clk_period;
		Addr <=  "00101010000101";
		Trees_din <= x"00092ad5";
		wait for Clk_period;
		Addr <=  "00101010000110";
		Trees_din <= x"ff922ad5";
		wait for Clk_period;
		Addr <=  "00101010000111";
		Trees_din <= x"0d004704";
		wait for Clk_period;
		Addr <=  "00101010001000";
		Trees_din <= x"ffcf2ad5";
		wait for Clk_period;
		Addr <=  "00101010001001";
		Trees_din <= x"00582ad5";
		wait for Clk_period;
		Addr <=  "00101010001010";
		Trees_din <= x"0007fa24";
		wait for Clk_period;
		Addr <=  "00101010001011";
		Trees_din <= x"1900a314";
		wait for Clk_period;
		Addr <=  "00101010001100";
		Trees_din <= x"14001804";
		wait for Clk_period;
		Addr <=  "00101010001101";
		Trees_din <= x"ffa42ad5";
		wait for Clk_period;
		Addr <=  "00101010001110";
		Trees_din <= x"06f24d08";
		wait for Clk_period;
		Addr <=  "00101010001111";
		Trees_din <= x"1d004604";
		wait for Clk_period;
		Addr <=  "00101010010000";
		Trees_din <= x"00592ad5";
		wait for Clk_period;
		Addr <=  "00101010010001";
		Trees_din <= x"ffd02ad5";
		wait for Clk_period;
		Addr <=  "00101010010010";
		Trees_din <= x"0bf94a04";
		wait for Clk_period;
		Addr <=  "00101010010011";
		Trees_din <= x"00212ad5";
		wait for Clk_period;
		Addr <=  "00101010010100";
		Trees_din <= x"00952ad5";
		wait for Clk_period;
		Addr <=  "00101010010101";
		Trees_din <= x"09005104";
		wait for Clk_period;
		Addr <=  "00101010010110";
		Trees_din <= x"00502ad5";
		wait for Clk_period;
		Addr <=  "00101010010111";
		Trees_din <= x"010ea204";
		wait for Clk_period;
		Addr <=  "00101010011000";
		Trees_din <= x"ff862ad5";
		wait for Clk_period;
		Addr <=  "00101010011001";
		Trees_din <= x"0ef9de04";
		wait for Clk_period;
		Addr <=  "00101010011010";
		Trees_din <= x"ffba2ad5";
		wait for Clk_period;
		Addr <=  "00101010011011";
		Trees_din <= x"002e2ad5";
		wait for Clk_period;
		Addr <=  "00101010011100";
		Trees_din <= x"1400c818";
		wait for Clk_period;
		Addr <=  "00101010011101";
		Trees_din <= x"11046d10";
		wait for Clk_period;
		Addr <=  "00101010011110";
		Trees_din <= x"0c021b08";
		wait for Clk_period;
		Addr <=  "00101010011111";
		Trees_din <= x"05f94a04";
		wait for Clk_period;
		Addr <=  "00101010100000";
		Trees_din <= x"ffff2ad5";
		wait for Clk_period;
		Addr <=  "00101010100001";
		Trees_din <= x"00662ad5";
		wait for Clk_period;
		Addr <=  "00101010100010";
		Trees_din <= x"07005a04";
		wait for Clk_period;
		Addr <=  "00101010100011";
		Trees_din <= x"ff8d2ad5";
		wait for Clk_period;
		Addr <=  "00101010100100";
		Trees_din <= x"00502ad5";
		wait for Clk_period;
		Addr <=  "00101010100101";
		Trees_din <= x"14008404";
		wait for Clk_period;
		Addr <=  "00101010100110";
		Trees_din <= x"ff8d2ad5";
		wait for Clk_period;
		Addr <=  "00101010100111";
		Trees_din <= x"00292ad5";
		wait for Clk_period;
		Addr <=  "00101010101000";
		Trees_din <= x"0d038c10";
		wait for Clk_period;
		Addr <=  "00101010101001";
		Trees_din <= x"0c033108";
		wait for Clk_period;
		Addr <=  "00101010101010";
		Trees_din <= x"06f66004";
		wait for Clk_period;
		Addr <=  "00101010101011";
		Trees_din <= x"ffdd2ad5";
		wait for Clk_period;
		Addr <=  "00101010101100";
		Trees_din <= x"00222ad5";
		wait for Clk_period;
		Addr <=  "00101010101101";
		Trees_din <= x"0bf94a04";
		wait for Clk_period;
		Addr <=  "00101010101110";
		Trees_din <= x"ffbc2ad5";
		wait for Clk_period;
		Addr <=  "00101010101111";
		Trees_din <= x"00532ad5";
		wait for Clk_period;
		Addr <=  "00101010110000";
		Trees_din <= x"03f30e04";
		wait for Clk_period;
		Addr <=  "00101010110001";
		Trees_din <= x"00502ad5";
		wait for Clk_period;
		Addr <=  "00101010110010";
		Trees_din <= x"14010404";
		wait for Clk_period;
		Addr <=  "00101010110011";
		Trees_din <= x"00192ad5";
		wait for Clk_period;
		Addr <=  "00101010110100";
		Trees_din <= x"ff7b2ad5";
		wait for Clk_period;
		Addr <=  "00101010110101";
		Trees_din <= x"0113e94c";
		wait for Clk_period;
		Addr <=  "00101010110110";
		Trees_din <= x"1e005b24";
		wait for Clk_period;
		Addr <=  "00101010110111";
		Trees_din <= x"0a04d620";
		wait for Clk_period;
		Addr <=  "00101010111000";
		Trees_din <= x"06f8b810";
		wait for Clk_period;
		Addr <=  "00101010111001";
		Trees_din <= x"06f71c08";
		wait for Clk_period;
		Addr <=  "00101010111010";
		Trees_din <= x"1f000004";
		wait for Clk_period;
		Addr <=  "00101010111011";
		Trees_din <= x"00232ba1";
		wait for Clk_period;
		Addr <=  "00101010111100";
		Trees_din <= x"ffbc2ba1";
		wait for Clk_period;
		Addr <=  "00101010111101";
		Trees_din <= x"0c021f04";
		wait for Clk_period;
		Addr <=  "00101010111110";
		Trees_din <= x"00872ba1";
		wait for Clk_period;
		Addr <=  "00101010111111";
		Trees_din <= x"00102ba1";
		wait for Clk_period;
		Addr <=  "00101011000000";
		Trees_din <= x"1e005708";
		wait for Clk_period;
		Addr <=  "00101011000001";
		Trees_din <= x"0200af04";
		wait for Clk_period;
		Addr <=  "00101011000010";
		Trees_din <= x"ffe02ba1";
		wait for Clk_period;
		Addr <=  "00101011000011";
		Trees_din <= x"ff892ba1";
		wait for Clk_period;
		Addr <=  "00101011000100";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00101011000101";
		Trees_din <= x"004f2ba1";
		wait for Clk_period;
		Addr <=  "00101011000110";
		Trees_din <= x"ffda2ba1";
		wait for Clk_period;
		Addr <=  "00101011000111";
		Trees_din <= x"ff8e2ba1";
		wait for Clk_period;
		Addr <=  "00101011001000";
		Trees_din <= x"1b003008";
		wait for Clk_period;
		Addr <=  "00101011001001";
		Trees_din <= x"0d020f04";
		wait for Clk_period;
		Addr <=  "00101011001010";
		Trees_din <= x"ffe72ba1";
		wait for Clk_period;
		Addr <=  "00101011001011";
		Trees_din <= x"ff6e2ba1";
		wait for Clk_period;
		Addr <=  "00101011001100";
		Trees_din <= x"1301ab10";
		wait for Clk_period;
		Addr <=  "00101011001101";
		Trees_din <= x"1203d308";
		wait for Clk_period;
		Addr <=  "00101011001110";
		Trees_din <= x"06f96104";
		wait for Clk_period;
		Addr <=  "00101011001111";
		Trees_din <= x"fff62ba1";
		wait for Clk_period;
		Addr <=  "00101011010000";
		Trees_din <= x"00262ba1";
		wait for Clk_period;
		Addr <=  "00101011010001";
		Trees_din <= x"07005204";
		wait for Clk_period;
		Addr <=  "00101011010010";
		Trees_din <= x"001c2ba1";
		wait for Clk_period;
		Addr <=  "00101011010011";
		Trees_din <= x"ff892ba1";
		wait for Clk_period;
		Addr <=  "00101011010100";
		Trees_din <= x"0bfb4c08";
		wait for Clk_period;
		Addr <=  "00101011010101";
		Trees_din <= x"10fbfc04";
		wait for Clk_period;
		Addr <=  "00101011010110";
		Trees_din <= x"00842ba1";
		wait for Clk_period;
		Addr <=  "00101011010111";
		Trees_din <= x"ffe02ba1";
		wait for Clk_period;
		Addr <=  "00101011011000";
		Trees_din <= x"0200c404";
		wait for Clk_period;
		Addr <=  "00101011011001";
		Trees_din <= x"00292ba1";
		wait for Clk_period;
		Addr <=  "00101011011010";
		Trees_din <= x"ff9b2ba1";
		wait for Clk_period;
		Addr <=  "00101011011011";
		Trees_din <= x"1a00e010";
		wait for Clk_period;
		Addr <=  "00101011011100";
		Trees_din <= x"1d004e08";
		wait for Clk_period;
		Addr <=  "00101011011101";
		Trees_din <= x"0015f004";
		wait for Clk_period;
		Addr <=  "00101011011110";
		Trees_din <= x"00792ba1";
		wait for Clk_period;
		Addr <=  "00101011011111";
		Trees_din <= x"00092ba1";
		wait for Clk_period;
		Addr <=  "00101011100000";
		Trees_din <= x"04f8eb04";
		wait for Clk_period;
		Addr <=  "00101011100001";
		Trees_din <= x"003d2ba1";
		wait for Clk_period;
		Addr <=  "00101011100010";
		Trees_din <= x"ffca2ba1";
		wait for Clk_period;
		Addr <=  "00101011100011";
		Trees_din <= x"1d003904";
		wait for Clk_period;
		Addr <=  "00101011100100";
		Trees_din <= x"00382ba1";
		wait for Clk_period;
		Addr <=  "00101011100101";
		Trees_din <= x"14020504";
		wait for Clk_period;
		Addr <=  "00101011100110";
		Trees_din <= x"fff02ba1";
		wait for Clk_period;
		Addr <=  "00101011100111";
		Trees_din <= x"ffb62ba1";
		wait for Clk_period;
		Addr <=  "00101011101000";
		Trees_din <= x"01114450";
		wait for Clk_period;
		Addr <=  "00101011101001";
		Trees_din <= x"03f78328";
		wait for Clk_period;
		Addr <=  "00101011101010";
		Trees_din <= x"03f63f14";
		wait for Clk_period;
		Addr <=  "00101011101011";
		Trees_din <= x"03f63510";
		wait for Clk_period;
		Addr <=  "00101011101100";
		Trees_din <= x"0d01af08";
		wait for Clk_period;
		Addr <=  "00101011101101";
		Trees_din <= x"06f76d04";
		wait for Clk_period;
		Addr <=  "00101011101110";
		Trees_din <= x"00322cbd";
		wait for Clk_period;
		Addr <=  "00101011101111";
		Trees_din <= x"ffbe2cbd";
		wait for Clk_period;
		Addr <=  "00101011110000";
		Trees_din <= x"03f30204";
		wait for Clk_period;
		Addr <=  "00101011110001";
		Trees_din <= x"00252cbd";
		wait for Clk_period;
		Addr <=  "00101011110010";
		Trees_din <= x"ff9d2cbd";
		wait for Clk_period;
		Addr <=  "00101011110011";
		Trees_din <= x"00872cbd";
		wait for Clk_period;
		Addr <=  "00101011110100";
		Trees_din <= x"0b04f20c";
		wait for Clk_period;
		Addr <=  "00101011110101";
		Trees_din <= x"02ff0b04";
		wait for Clk_period;
		Addr <=  "00101011110110";
		Trees_din <= x"00392cbd";
		wait for Clk_period;
		Addr <=  "00101011110111";
		Trees_din <= x"0a02f104";
		wait for Clk_period;
		Addr <=  "00101011111000";
		Trees_din <= x"ff7d2cbd";
		wait for Clk_period;
		Addr <=  "00101011111001";
		Trees_din <= x"fffa2cbd";
		wait for Clk_period;
		Addr <=  "00101011111010";
		Trees_din <= x"06f3a804";
		wait for Clk_period;
		Addr <=  "00101011111011";
		Trees_din <= x"005a2cbd";
		wait for Clk_period;
		Addr <=  "00101011111100";
		Trees_din <= x"ffda2cbd";
		wait for Clk_period;
		Addr <=  "00101011111101";
		Trees_din <= x"01107320";
		wait for Clk_period;
		Addr <=  "00101011111110";
		Trees_din <= x"0b049410";
		wait for Clk_period;
		Addr <=  "00101011111111";
		Trees_din <= x"0b046408";
		wait for Clk_period;
		Addr <=  "00101100000000";
		Trees_din <= x"05fda304";
		wait for Clk_period;
		Addr <=  "00101100000001";
		Trees_din <= x"00082cbd";
		wait for Clk_period;
		Addr <=  "00101100000010";
		Trees_din <= x"ffc92cbd";
		wait for Clk_period;
		Addr <=  "00101100000011";
		Trees_din <= x"0d032504";
		wait for Clk_period;
		Addr <=  "00101100000100";
		Trees_din <= x"00882cbd";
		wait for Clk_period;
		Addr <=  "00101100000101";
		Trees_din <= x"fff12cbd";
		wait for Clk_period;
		Addr <=  "00101100000110";
		Trees_din <= x"09005908";
		wait for Clk_period;
		Addr <=  "00101100000111";
		Trees_din <= x"15009904";
		wait for Clk_period;
		Addr <=  "00101100001000";
		Trees_din <= x"00282cbd";
		wait for Clk_period;
		Addr <=  "00101100001001";
		Trees_din <= x"ffcd2cbd";
		wait for Clk_period;
		Addr <=  "00101100001010";
		Trees_din <= x"0efdd204";
		wait for Clk_period;
		Addr <=  "00101100001011";
		Trees_din <= x"000f2cbd";
		wait for Clk_period;
		Addr <=  "00101100001100";
		Trees_din <= x"ff6e2cbd";
		wait for Clk_period;
		Addr <=  "00101100001101";
		Trees_din <= x"1b003604";
		wait for Clk_period;
		Addr <=  "00101100001110";
		Trees_din <= x"001c2cbd";
		wait for Clk_period;
		Addr <=  "00101100001111";
		Trees_din <= x"00792cbd";
		wait for Clk_period;
		Addr <=  "00101100010000";
		Trees_din <= x"0b049930";
		wait for Clk_period;
		Addr <=  "00101100010001";
		Trees_din <= x"0b027d14";
		wait for Clk_period;
		Addr <=  "00101100010010";
		Trees_din <= x"0f000104";
		wait for Clk_period;
		Addr <=  "00101100010011";
		Trees_din <= x"ffad2cbd";
		wait for Clk_period;
		Addr <=  "00101100010100";
		Trees_din <= x"00126b08";
		wait for Clk_period;
		Addr <=  "00101100010101";
		Trees_din <= x"0d03a504";
		wait for Clk_period;
		Addr <=  "00101100010110";
		Trees_din <= x"00672cbd";
		wait for Clk_period;
		Addr <=  "00101100010111";
		Trees_din <= x"fff42cbd";
		wait for Clk_period;
		Addr <=  "00101100011000";
		Trees_din <= x"15009304";
		wait for Clk_period;
		Addr <=  "00101100011001";
		Trees_din <= x"ffb52cbd";
		wait for Clk_period;
		Addr <=  "00101100011010";
		Trees_din <= x"00232cbd";
		wait for Clk_period;
		Addr <=  "00101100011011";
		Trees_din <= x"1401770c";
		wait for Clk_period;
		Addr <=  "00101100011100";
		Trees_din <= x"03f82f08";
		wait for Clk_period;
		Addr <=  "00101100011101";
		Trees_din <= x"1a00bc04";
		wait for Clk_period;
		Addr <=  "00101100011110";
		Trees_din <= x"fffd2cbd";
		wait for Clk_period;
		Addr <=  "00101100011111";
		Trees_din <= x"006b2cbd";
		wait for Clk_period;
		Addr <=  "00101100100000";
		Trees_din <= x"ffcd2cbd";
		wait for Clk_period;
		Addr <=  "00101100100001";
		Trees_din <= x"000c5808";
		wait for Clk_period;
		Addr <=  "00101100100010";
		Trees_din <= x"13f9c904";
		wait for Clk_period;
		Addr <=  "00101100100011";
		Trees_din <= x"ffda2cbd";
		wait for Clk_period;
		Addr <=  "00101100100100";
		Trees_din <= x"00592cbd";
		wait for Clk_period;
		Addr <=  "00101100100101";
		Trees_din <= x"0802c204";
		wait for Clk_period;
		Addr <=  "00101100100110";
		Trees_din <= x"ff6c2cbd";
		wait for Clk_period;
		Addr <=  "00101100100111";
		Trees_din <= x"fffa2cbd";
		wait for Clk_period;
		Addr <=  "00101100101000";
		Trees_din <= x"1500a208";
		wait for Clk_period;
		Addr <=  "00101100101001";
		Trees_din <= x"00148704";
		wait for Clk_period;
		Addr <=  "00101100101010";
		Trees_din <= x"00822cbd";
		wait for Clk_period;
		Addr <=  "00101100101011";
		Trees_din <= x"00132cbd";
		wait for Clk_period;
		Addr <=  "00101100101100";
		Trees_din <= x"12001904";
		wait for Clk_period;
		Addr <=  "00101100101101";
		Trees_din <= x"ffe22cbd";
		wait for Clk_period;
		Addr <=  "00101100101110";
		Trees_din <= x"000a2cbd";
		wait for Clk_period;
		Addr <=  "00101100101111";
		Trees_din <= x"0105aa34";
		wait for Clk_period;
		Addr <=  "00101100110000";
		Trees_din <= x"03fc9708";
		wait for Clk_period;
		Addr <=  "00101100110001";
		Trees_din <= x"0c006e04";
		wait for Clk_period;
		Addr <=  "00101100110010";
		Trees_din <= x"001d2df1";
		wait for Clk_period;
		Addr <=  "00101100110011";
		Trees_din <= x"ff7d2df1";
		wait for Clk_period;
		Addr <=  "00101100110100";
		Trees_din <= x"04025d14";
		wait for Clk_period;
		Addr <=  "00101100110101";
		Trees_din <= x"14005204";
		wait for Clk_period;
		Addr <=  "00101100110110";
		Trees_din <= x"ffa42df1";
		wait for Clk_period;
		Addr <=  "00101100110111";
		Trees_din <= x"08019908";
		wait for Clk_period;
		Addr <=  "00101100111000";
		Trees_din <= x"19009104";
		wait for Clk_period;
		Addr <=  "00101100111001";
		Trees_din <= x"fff92df1";
		wait for Clk_period;
		Addr <=  "00101100111010";
		Trees_din <= x"00672df1";
		wait for Clk_period;
		Addr <=  "00101100111011";
		Trees_din <= x"08030104";
		wait for Clk_period;
		Addr <=  "00101100111100";
		Trees_din <= x"ff912df1";
		wait for Clk_period;
		Addr <=  "00101100111101";
		Trees_din <= x"00312df1";
		wait for Clk_period;
		Addr <=  "00101100111110";
		Trees_din <= x"0f000f08";
		wait for Clk_period;
		Addr <=  "00101100111111";
		Trees_din <= x"1900a104";
		wait for Clk_period;
		Addr <=  "00101101000000";
		Trees_din <= x"fffb2df1";
		wait for Clk_period;
		Addr <=  "00101101000001";
		Trees_din <= x"00682df1";
		wait for Clk_period;
		Addr <=  "00101101000010";
		Trees_din <= x"0f01d108";
		wait for Clk_period;
		Addr <=  "00101101000011";
		Trees_din <= x"16017504";
		wait for Clk_period;
		Addr <=  "00101101000100";
		Trees_din <= x"ffe42df1";
		wait for Clk_period;
		Addr <=  "00101101000101";
		Trees_din <= x"ff7b2df1";
		wait for Clk_period;
		Addr <=  "00101101000110";
		Trees_din <= x"17000004";
		wait for Clk_period;
		Addr <=  "00101101000111";
		Trees_din <= x"ff9c2df1";
		wait for Clk_period;
		Addr <=  "00101101001000";
		Trees_din <= x"00162df1";
		wait for Clk_period;
		Addr <=  "00101101001001";
		Trees_din <= x"0f003e30";
		wait for Clk_period;
		Addr <=  "00101101001010";
		Trees_din <= x"0f001f1c";
		wait for Clk_period;
		Addr <=  "00101101001011";
		Trees_din <= x"1700150c";
		wait for Clk_period;
		Addr <=  "00101101001100";
		Trees_din <= x"1500a008";
		wait for Clk_period;
		Addr <=  "00101101001101";
		Trees_din <= x"01081404";
		wait for Clk_period;
		Addr <=  "00101101001110";
		Trees_din <= x"fff82df1";
		wait for Clk_period;
		Addr <=  "00101101001111";
		Trees_din <= x"00712df1";
		wait for Clk_period;
		Addr <=  "00101101010000";
		Trees_din <= x"ffdb2df1";
		wait for Clk_period;
		Addr <=  "00101101010001";
		Trees_din <= x"0e009508";
		wait for Clk_period;
		Addr <=  "00101101010010";
		Trees_din <= x"09005a04";
		wait for Clk_period;
		Addr <=  "00101101010011";
		Trees_din <= x"002f2df1";
		wait for Clk_period;
		Addr <=  "00101101010100";
		Trees_din <= x"ff982df1";
		wait for Clk_period;
		Addr <=  "00101101010101";
		Trees_din <= x"0f001404";
		wait for Clk_period;
		Addr <=  "00101101010110";
		Trees_din <= x"ffb22df1";
		wait for Clk_period;
		Addr <=  "00101101010111";
		Trees_din <= x"00272df1";
		wait for Clk_period;
		Addr <=  "00101101011000";
		Trees_din <= x"01114410";
		wait for Clk_period;
		Addr <=  "00101101011001";
		Trees_din <= x"1d003b08";
		wait for Clk_period;
		Addr <=  "00101101011010";
		Trees_din <= x"14007804";
		wait for Clk_period;
		Addr <=  "00101101011011";
		Trees_din <= x"004a2df1";
		wait for Clk_period;
		Addr <=  "00101101011100";
		Trees_din <= x"ffc52df1";
		wait for Clk_period;
		Addr <=  "00101101011101";
		Trees_din <= x"0af77a04";
		wait for Clk_period;
		Addr <=  "00101101011110";
		Trees_din <= x"00062df1";
		wait for Clk_period;
		Addr <=  "00101101011111";
		Trees_din <= x"ff792df1";
		wait for Clk_period;
		Addr <=  "00101101100000";
		Trees_din <= x"00462df1";
		wait for Clk_period;
		Addr <=  "00101101100001";
		Trees_din <= x"0200e118";
		wait for Clk_period;
		Addr <=  "00101101100010";
		Trees_din <= x"16000308";
		wait for Clk_period;
		Addr <=  "00101101100011";
		Trees_din <= x"02002404";
		wait for Clk_period;
		Addr <=  "00101101100100";
		Trees_din <= x"ffa02df1";
		wait for Clk_period;
		Addr <=  "00101101100101";
		Trees_din <= x"000e2df1";
		wait for Clk_period;
		Addr <=  "00101101100110";
		Trees_din <= x"09005a08";
		wait for Clk_period;
		Addr <=  "00101101100111";
		Trees_din <= x"16039604";
		wait for Clk_period;
		Addr <=  "00101101101000";
		Trees_din <= x"00142df1";
		wait for Clk_period;
		Addr <=  "00101101101001";
		Trees_din <= x"00652df1";
		wait for Clk_period;
		Addr <=  "00101101101010";
		Trees_din <= x"0f013204";
		wait for Clk_period;
		Addr <=  "00101101101011";
		Trees_din <= x"fff22df1";
		wait for Clk_period;
		Addr <=  "00101101101100";
		Trees_din <= x"008d2df1";
		wait for Clk_period;
		Addr <=  "00101101101101";
		Trees_din <= x"02019d10";
		wait for Clk_period;
		Addr <=  "00101101101110";
		Trees_din <= x"06f7d008";
		wait for Clk_period;
		Addr <=  "00101101101111";
		Trees_din <= x"06f23704";
		wait for Clk_period;
		Addr <=  "00101101110000";
		Trees_din <= x"002c2df1";
		wait for Clk_period;
		Addr <=  "00101101110001";
		Trees_din <= x"ff892df1";
		wait for Clk_period;
		Addr <=  "00101101110010";
		Trees_din <= x"1602fa04";
		wait for Clk_period;
		Addr <=  "00101101110011";
		Trees_din <= x"ffe12df1";
		wait for Clk_period;
		Addr <=  "00101101110100";
		Trees_din <= x"00852df1";
		wait for Clk_period;
		Addr <=  "00101101110101";
		Trees_din <= x"13fa0b08";
		wait for Clk_period;
		Addr <=  "00101101110110";
		Trees_din <= x"03f93a04";
		wait for Clk_period;
		Addr <=  "00101101110111";
		Trees_din <= x"00122df1";
		wait for Clk_period;
		Addr <=  "00101101111000";
		Trees_din <= x"ffb62df1";
		wait for Clk_period;
		Addr <=  "00101101111001";
		Trees_din <= x"08018d04";
		wait for Clk_period;
		Addr <=  "00101101111010";
		Trees_din <= x"ffff2df1";
		wait for Clk_period;
		Addr <=  "00101101111011";
		Trees_din <= x"00332df1";
		wait for Clk_period;
		Addr <=  "00101101111100";
		Trees_din <= x"0105aa34";
		wait for Clk_period;
		Addr <=  "00101101111101";
		Trees_din <= x"03fc9708";
		wait for Clk_period;
		Addr <=  "00101101111110";
		Trees_din <= x"0c006e04";
		wait for Clk_period;
		Addr <=  "00101101111111";
		Trees_din <= x"00172ed5";
		wait for Clk_period;
		Addr <=  "00101110000000";
		Trees_din <= x"ff802ed5";
		wait for Clk_period;
		Addr <=  "00101110000001";
		Trees_din <= x"04025d14";
		wait for Clk_period;
		Addr <=  "00101110000010";
		Trees_din <= x"14005204";
		wait for Clk_period;
		Addr <=  "00101110000011";
		Trees_din <= x"ffa82ed5";
		wait for Clk_period;
		Addr <=  "00101110000100";
		Trees_din <= x"0c016e08";
		wait for Clk_period;
		Addr <=  "00101110000101";
		Trees_din <= x"19009104";
		wait for Clk_period;
		Addr <=  "00101110000110";
		Trees_din <= x"ffd32ed5";
		wait for Clk_period;
		Addr <=  "00101110000111";
		Trees_din <= x"00732ed5";
		wait for Clk_period;
		Addr <=  "00101110001000";
		Trees_din <= x"00090504";
		wait for Clk_period;
		Addr <=  "00101110001001";
		Trees_din <= x"00232ed5";
		wait for Clk_period;
		Addr <=  "00101110001010";
		Trees_din <= x"ffb42ed5";
		wait for Clk_period;
		Addr <=  "00101110001011";
		Trees_din <= x"0f000f08";
		wait for Clk_period;
		Addr <=  "00101110001100";
		Trees_din <= x"1900a104";
		wait for Clk_period;
		Addr <=  "00101110001101";
		Trees_din <= x"fff92ed5";
		wait for Clk_period;
		Addr <=  "00101110001110";
		Trees_din <= x"005d2ed5";
		wait for Clk_period;
		Addr <=  "00101110001111";
		Trees_din <= x"12025208";
		wait for Clk_period;
		Addr <=  "00101110010000";
		Trees_din <= x"1a009c04";
		wait for Clk_period;
		Addr <=  "00101110010001";
		Trees_din <= x"fffa2ed5";
		wait for Clk_period;
		Addr <=  "00101110010010";
		Trees_din <= x"ff7c2ed5";
		wait for Clk_period;
		Addr <=  "00101110010011";
		Trees_din <= x"0bfa8104";
		wait for Clk_period;
		Addr <=  "00101110010100";
		Trees_din <= x"003a2ed5";
		wait for Clk_period;
		Addr <=  "00101110010101";
		Trees_din <= x"ffb22ed5";
		wait for Clk_period;
		Addr <=  "00101110010110";
		Trees_din <= x"0bf95618";
		wait for Clk_period;
		Addr <=  "00101110010111";
		Trees_din <= x"09005710";
		wait for Clk_period;
		Addr <=  "00101110011000";
		Trees_din <= x"1603e80c";
		wait for Clk_period;
		Addr <=  "00101110011001";
		Trees_din <= x"10055408";
		wait for Clk_period;
		Addr <=  "00101110011010";
		Trees_din <= x"0207bf04";
		wait for Clk_period;
		Addr <=  "00101110011011";
		Trees_din <= x"00492ed5";
		wait for Clk_period;
		Addr <=  "00101110011100";
		Trees_din <= x"ffe12ed5";
		wait for Clk_period;
		Addr <=  "00101110011101";
		Trees_din <= x"ffb22ed5";
		wait for Clk_period;
		Addr <=  "00101110011110";
		Trees_din <= x"ffa72ed5";
		wait for Clk_period;
		Addr <=  "00101110011111";
		Trees_din <= x"1a00ca04";
		wait for Clk_period;
		Addr <=  "00101110100000";
		Trees_din <= x"ff872ed5";
		wait for Clk_period;
		Addr <=  "00101110100001";
		Trees_din <= x"ffeb2ed5";
		wait for Clk_period;
		Addr <=  "00101110100010";
		Trees_din <= x"0d03ea20";
		wait for Clk_period;
		Addr <=  "00101110100011";
		Trees_din <= x"1c003210";
		wait for Clk_period;
		Addr <=  "00101110100100";
		Trees_din <= x"1e005b08";
		wait for Clk_period;
		Addr <=  "00101110100101";
		Trees_din <= x"13019204";
		wait for Clk_period;
		Addr <=  "00101110100110";
		Trees_din <= x"00212ed5";
		wait for Clk_period;
		Addr <=  "00101110100111";
		Trees_din <= x"ffa72ed5";
		wait for Clk_period;
		Addr <=  "00101110101000";
		Trees_din <= x"1201f904";
		wait for Clk_period;
		Addr <=  "00101110101001";
		Trees_din <= x"00022ed5";
		wait for Clk_period;
		Addr <=  "00101110101010";
		Trees_din <= x"ffae2ed5";
		wait for Clk_period;
		Addr <=  "00101110101011";
		Trees_din <= x"0bf97c08";
		wait for Clk_period;
		Addr <=  "00101110101100";
		Trees_din <= x"09005504";
		wait for Clk_period;
		Addr <=  "00101110101101";
		Trees_din <= x"ffec2ed5";
		wait for Clk_period;
		Addr <=  "00101110101110";
		Trees_din <= x"00852ed5";
		wait for Clk_period;
		Addr <=  "00101110101111";
		Trees_din <= x"06f4cb04";
		wait for Clk_period;
		Addr <=  "00101110110000";
		Trees_din <= x"00232ed5";
		wait for Clk_period;
		Addr <=  "00101110110001";
		Trees_din <= x"fff92ed5";
		wait for Clk_period;
		Addr <=  "00101110110010";
		Trees_din <= x"07005a04";
		wait for Clk_period;
		Addr <=  "00101110110011";
		Trees_din <= x"ff9d2ed5";
		wait for Clk_period;
		Addr <=  "00101110110100";
		Trees_din <= x"fff72ed5";
		wait for Clk_period;
		Addr <=  "00101110110101";
		Trees_din <= x"010d4f40";
		wait for Clk_period;
		Addr <=  "00101110110110";
		Trees_din <= x"13014d1c";
		wait for Clk_period;
		Addr <=  "00101110110111";
		Trees_din <= x"13013a18";
		wait for Clk_period;
		Addr <=  "00101110111000";
		Trees_din <= x"03f6f40c";
		wait for Clk_period;
		Addr <=  "00101110111001";
		Trees_din <= x"10028708";
		wait for Clk_period;
		Addr <=  "00101110111010";
		Trees_din <= x"04f80404";
		wait for Clk_period;
		Addr <=  "00101110111011";
		Trees_din <= x"ffbe3009";
		wait for Clk_period;
		Addr <=  "00101110111100";
		Trees_din <= x"00463009";
		wait for Clk_period;
		Addr <=  "00101110111101";
		Trees_din <= x"ff883009";
		wait for Clk_period;
		Addr <=  "00101110111110";
		Trees_din <= x"010d2808";
		wait for Clk_period;
		Addr <=  "00101110111111";
		Trees_din <= x"010cb404";
		wait for Clk_period;
		Addr <=  "00101111000000";
		Trees_din <= x"ffff3009";
		wait for Clk_period;
		Addr <=  "00101111000001";
		Trees_din <= x"00423009";
		wait for Clk_period;
		Addr <=  "00101111000010";
		Trees_din <= x"ffa23009";
		wait for Clk_period;
		Addr <=  "00101111000011";
		Trees_din <= x"00753009";
		wait for Clk_period;
		Addr <=  "00101111000100";
		Trees_din <= x"06f3580c";
		wait for Clk_period;
		Addr <=  "00101111000101";
		Trees_din <= x"1401dd04";
		wait for Clk_period;
		Addr <=  "00101111000110";
		Trees_din <= x"ffd33009";
		wait for Clk_period;
		Addr <=  "00101111000111";
		Trees_din <= x"07005704";
		wait for Clk_period;
		Addr <=  "00101111001000";
		Trees_din <= x"00253009";
		wait for Clk_period;
		Addr <=  "00101111001001";
		Trees_din <= x"00783009";
		wait for Clk_period;
		Addr <=  "00101111001010";
		Trees_din <= x"0d037310";
		wait for Clk_period;
		Addr <=  "00101111001011";
		Trees_din <= x"0e035208";
		wait for Clk_period;
		Addr <=  "00101111001100";
		Trees_din <= x"03fc1504";
		wait for Clk_period;
		Addr <=  "00101111001101";
		Trees_din <= x"ffac3009";
		wait for Clk_period;
		Addr <=  "00101111001110";
		Trees_din <= x"00213009";
		wait for Clk_period;
		Addr <=  "00101111001111";
		Trees_din <= x"09005804";
		wait for Clk_period;
		Addr <=  "00101111010000";
		Trees_din <= x"ff6d3009";
		wait for Clk_period;
		Addr <=  "00101111010001";
		Trees_din <= x"ffc93009";
		wait for Clk_period;
		Addr <=  "00101111010010";
		Trees_din <= x"01090e04";
		wait for Clk_period;
		Addr <=  "00101111010011";
		Trees_din <= x"ffd33009";
		wait for Clk_period;
		Addr <=  "00101111010100";
		Trees_din <= x"004c3009";
		wait for Clk_period;
		Addr <=  "00101111010101";
		Trees_din <= x"03f9b834";
		wait for Clk_period;
		Addr <=  "00101111010110";
		Trees_din <= x"1403ab20";
		wait for Clk_period;
		Addr <=  "00101111010111";
		Trees_din <= x"1400c810";
		wait for Clk_period;
		Addr <=  "00101111011000";
		Trees_din <= x"11046d08";
		wait for Clk_period;
		Addr <=  "00101111011001";
		Trees_din <= x"0012ed04";
		wait for Clk_period;
		Addr <=  "00101111011010";
		Trees_din <= x"00403009";
		wait for Clk_period;
		Addr <=  "00101111011011";
		Trees_din <= x"ffdf3009";
		wait for Clk_period;
		Addr <=  "00101111011100";
		Trees_din <= x"0801d404";
		wait for Clk_period;
		Addr <=  "00101111011101";
		Trees_din <= x"ffa33009";
		wait for Clk_period;
		Addr <=  "00101111011110";
		Trees_din <= x"00083009";
		wait for Clk_period;
		Addr <=  "00101111011111";
		Trees_din <= x"05f9bd08";
		wait for Clk_period;
		Addr <=  "00101111100000";
		Trees_din <= x"0c028604";
		wait for Clk_period;
		Addr <=  "00101111100001";
		Trees_din <= x"ffd53009";
		wait for Clk_period;
		Addr <=  "00101111100010";
		Trees_din <= x"003b3009";
		wait for Clk_period;
		Addr <=  "00101111100011";
		Trees_din <= x"05fa8c04";
		wait for Clk_period;
		Addr <=  "00101111100100";
		Trees_din <= x"ff9b3009";
		wait for Clk_period;
		Addr <=  "00101111100101";
		Trees_din <= x"fff43009";
		wait for Clk_period;
		Addr <=  "00101111100110";
		Trees_din <= x"10fade04";
		wait for Clk_period;
		Addr <=  "00101111100111";
		Trees_din <= x"ffc33009";
		wait for Clk_period;
		Addr <=  "00101111101000";
		Trees_din <= x"12ff1908";
		wait for Clk_period;
		Addr <=  "00101111101001";
		Trees_din <= x"03f74704";
		wait for Clk_period;
		Addr <=  "00101111101010";
		Trees_din <= x"ffbb3009";
		wait for Clk_period;
		Addr <=  "00101111101011";
		Trees_din <= x"002a3009";
		wait for Clk_period;
		Addr <=  "00101111101100";
		Trees_din <= x"03f4a004";
		wait for Clk_period;
		Addr <=  "00101111101101";
		Trees_din <= x"00113009";
		wait for Clk_period;
		Addr <=  "00101111101110";
		Trees_din <= x"007e3009";
		wait for Clk_period;
		Addr <=  "00101111101111";
		Trees_din <= x"13fdb118";
		wait for Clk_period;
		Addr <=  "00101111110000";
		Trees_din <= x"10040610";
		wait for Clk_period;
		Addr <=  "00101111110001";
		Trees_din <= x"17000408";
		wait for Clk_period;
		Addr <=  "00101111110010";
		Trees_din <= x"14037804";
		wait for Clk_period;
		Addr <=  "00101111110011";
		Trees_din <= x"005c3009";
		wait for Clk_period;
		Addr <=  "00101111110100";
		Trees_din <= x"ffc43009";
		wait for Clk_period;
		Addr <=  "00101111110101";
		Trees_din <= x"15009c04";
		wait for Clk_period;
		Addr <=  "00101111110110";
		Trees_din <= x"ffe23009";
		wait for Clk_period;
		Addr <=  "00101111110111";
		Trees_din <= x"ff773009";
		wait for Clk_period;
		Addr <=  "00101111111000";
		Trees_din <= x"08009604";
		wait for Clk_period;
		Addr <=  "00101111111001";
		Trees_din <= x"00083009";
		wait for Clk_period;
		Addr <=  "00101111111010";
		Trees_din <= x"006a3009";
		wait for Clk_period;
		Addr <=  "00101111111011";
		Trees_din <= x"0f000604";
		wait for Clk_period;
		Addr <=  "00101111111100";
		Trees_din <= x"ffda3009";
		wait for Clk_period;
		Addr <=  "00101111111101";
		Trees_din <= x"00fd6404";
		wait for Clk_period;
		Addr <=  "00101111111110";
		Trees_din <= x"ffe83009";
		wait for Clk_period;
		Addr <=  "00101111111111";
		Trees_din <= x"0d035b04";
		wait for Clk_period;
		Addr <=  "00110000000000";
		Trees_din <= x"00893009";
		wait for Clk_period;
		Addr <=  "00110000000001";
		Trees_din <= x"002d3009";
		wait for Clk_period;
		Addr <=  "00110000000010";
		Trees_din <= x"01164234";
		wait for Clk_period;
		Addr <=  "00110000000011";
		Trees_din <= x"1303b428";
		wait for Clk_period;
		Addr <=  "00110000000100";
		Trees_din <= x"0101750c";
		wait for Clk_period;
		Addr <=  "00110000000101";
		Trees_din <= x"02026c04";
		wait for Clk_period;
		Addr <=  "00110000000110";
		Trees_din <= x"ff91307d";
		wait for Clk_period;
		Addr <=  "00110000000111";
		Trees_din <= x"0203f904";
		wait for Clk_period;
		Addr <=  "00110000001000";
		Trees_din <= x"0049307d";
		wait for Clk_period;
		Addr <=  "00110000001001";
		Trees_din <= x"ffc4307d";
		wait for Clk_period;
		Addr <=  "00110000001010";
		Trees_din <= x"1500af10";
		wait for Clk_period;
		Addr <=  "00110000001011";
		Trees_din <= x"1b002908";
		wait for Clk_period;
		Addr <=  "00110000001100";
		Trees_din <= x"0f017304";
		wait for Clk_period;
		Addr <=  "00110000001101";
		Trees_din <= x"ff86307d";
		wait for Clk_period;
		Addr <=  "00110000001110";
		Trees_din <= x"000c307d";
		wait for Clk_period;
		Addr <=  "00110000001111";
		Trees_din <= x"07004c04";
		wait for Clk_period;
		Addr <=  "00110000010000";
		Trees_din <= x"0028307d";
		wait for Clk_period;
		Addr <=  "00110000010001";
		Trees_din <= x"fffd307d";
		wait for Clk_period;
		Addr <=  "00110000010010";
		Trees_din <= x"07004e04";
		wait for Clk_period;
		Addr <=  "00110000010011";
		Trees_din <= x"ffc4307d";
		wait for Clk_period;
		Addr <=  "00110000010100";
		Trees_din <= x"1e004d04";
		wait for Clk_period;
		Addr <=  "00110000010101";
		Trees_din <= x"007b307d";
		wait for Clk_period;
		Addr <=  "00110000010110";
		Trees_din <= x"0001307d";
		wait for Clk_period;
		Addr <=  "00110000010111";
		Trees_din <= x"10fc3608";
		wait for Clk_period;
		Addr <=  "00110000011000";
		Trees_din <= x"18003f04";
		wait for Clk_period;
		Addr <=  "00110000011001";
		Trees_din <= x"006e307d";
		wait for Clk_period;
		Addr <=  "00110000011010";
		Trees_din <= x"0018307d";
		wait for Clk_period;
		Addr <=  "00110000011011";
		Trees_din <= x"ffec307d";
		wait for Clk_period;
		Addr <=  "00110000011100";
		Trees_din <= x"08008a04";
		wait for Clk_period;
		Addr <=  "00110000011101";
		Trees_din <= x"000b307d";
		wait for Clk_period;
		Addr <=  "00110000011110";
		Trees_din <= x"0056307d";
		wait for Clk_period;
		Addr <=  "00110000011111";
		Trees_din <= x"010a1f48";
		wait for Clk_period;
		Addr <=  "00110000100000";
		Trees_din <= x"09005620";
		wait for Clk_period;
		Addr <=  "00110000100001";
		Trees_din <= x"04f88108";
		wait for Clk_period;
		Addr <=  "00110000100010";
		Trees_din <= x"0a043904";
		wait for Clk_period;
		Addr <=  "00110000100011";
		Trees_din <= x"ff8431b9";
		wait for Clk_period;
		Addr <=  "00110000100100";
		Trees_din <= x"002a31b9";
		wait for Clk_period;
		Addr <=  "00110000100101";
		Trees_din <= x"04f94b08";
		wait for Clk_period;
		Addr <=  "00110000100110";
		Trees_din <= x"0f01b404";
		wait for Clk_period;
		Addr <=  "00110000100111";
		Trees_din <= x"ffd531b9";
		wait for Clk_period;
		Addr <=  "00110000101000";
		Trees_din <= x"007831b9";
		wait for Clk_period;
		Addr <=  "00110000101001";
		Trees_din <= x"020b0108";
		wait for Clk_period;
		Addr <=  "00110000101010";
		Trees_din <= x"1a00e204";
		wait for Clk_period;
		Addr <=  "00110000101011";
		Trees_din <= x"ffc631b9";
		wait for Clk_period;
		Addr <=  "00110000101100";
		Trees_din <= x"000b31b9";
		wait for Clk_period;
		Addr <=  "00110000101101";
		Trees_din <= x"00042104";
		wait for Clk_period;
		Addr <=  "00110000101110";
		Trees_din <= x"ffca31b9";
		wait for Clk_period;
		Addr <=  "00110000101111";
		Trees_din <= x"005931b9";
		wait for Clk_period;
		Addr <=  "00110000110000";
		Trees_din <= x"04fd7914";
		wait for Clk_period;
		Addr <=  "00110000110001";
		Trees_din <= x"1e006304";
		wait for Clk_period;
		Addr <=  "00110000110010";
		Trees_din <= x"ffb731b9";
		wait for Clk_period;
		Addr <=  "00110000110011";
		Trees_din <= x"1e007808";
		wait for Clk_period;
		Addr <=  "00110000110100";
		Trees_din <= x"05fbfd04";
		wait for Clk_period;
		Addr <=  "00110000110101";
		Trees_din <= x"008031b9";
		wait for Clk_period;
		Addr <=  "00110000110110";
		Trees_din <= x"000231b9";
		wait for Clk_period;
		Addr <=  "00110000110111";
		Trees_din <= x"0008bf04";
		wait for Clk_period;
		Addr <=  "00110000111000";
		Trees_din <= x"004031b9";
		wait for Clk_period;
		Addr <=  "00110000111001";
		Trees_din <= x"ff9331b9";
		wait for Clk_period;
		Addr <=  "00110000111010";
		Trees_din <= x"03fbf604";
		wait for Clk_period;
		Addr <=  "00110000111011";
		Trees_din <= x"ff8831b9";
		wait for Clk_period;
		Addr <=  "00110000111100";
		Trees_din <= x"0bf9bc08";
		wait for Clk_period;
		Addr <=  "00110000111101";
		Trees_din <= x"1c003b04";
		wait for Clk_period;
		Addr <=  "00110000111110";
		Trees_din <= x"ff8431b9";
		wait for Clk_period;
		Addr <=  "00110000111111";
		Trees_din <= x"000f31b9";
		wait for Clk_period;
		Addr <=  "00110001000000";
		Trees_din <= x"0f000b04";
		wait for Clk_period;
		Addr <=  "00110001000001";
		Trees_din <= x"ffa331b9";
		wait for Clk_period;
		Addr <=  "00110001000010";
		Trees_din <= x"002731b9";
		wait for Clk_period;
		Addr <=  "00110001000011";
		Trees_din <= x"0007fa2c";
		wait for Clk_period;
		Addr <=  "00110001000100";
		Trees_din <= x"1900a118";
		wait for Clk_period;
		Addr <=  "00110001000101";
		Trees_din <= x"07005c10";
		wait for Clk_period;
		Addr <=  "00110001000110";
		Trees_din <= x"00fde508";
		wait for Clk_period;
		Addr <=  "00110001000111";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00110001001000";
		Trees_din <= x"003731b9";
		wait for Clk_period;
		Addr <=  "00110001001001";
		Trees_din <= x"ffb231b9";
		wait for Clk_period;
		Addr <=  "00110001001010";
		Trees_din <= x"15007c04";
		wait for Clk_period;
		Addr <=  "00110001001011";
		Trees_din <= x"ffe931b9";
		wait for Clk_period;
		Addr <=  "00110001001100";
		Trees_din <= x"007631b9";
		wait for Clk_period;
		Addr <=  "00110001001101";
		Trees_din <= x"06f52a04";
		wait for Clk_period;
		Addr <=  "00110001001110";
		Trees_din <= x"ffac31b9";
		wait for Clk_period;
		Addr <=  "00110001001111";
		Trees_din <= x"002c31b9";
		wait for Clk_period;
		Addr <=  "00110001010000";
		Trees_din <= x"09005004";
		wait for Clk_period;
		Addr <=  "00110001010001";
		Trees_din <= x"006a31b9";
		wait for Clk_period;
		Addr <=  "00110001010010";
		Trees_din <= x"0202a008";
		wait for Clk_period;
		Addr <=  "00110001010011";
		Trees_din <= x"04065f04";
		wait for Clk_period;
		Addr <=  "00110001010100";
		Trees_din <= x"006131b9";
		wait for Clk_period;
		Addr <=  "00110001010101";
		Trees_din <= x"ffc331b9";
		wait for Clk_period;
		Addr <=  "00110001010110";
		Trees_din <= x"010ea204";
		wait for Clk_period;
		Addr <=  "00110001010111";
		Trees_din <= x"ff7a31b9";
		wait for Clk_period;
		Addr <=  "00110001011000";
		Trees_din <= x"000431b9";
		wait for Clk_period;
		Addr <=  "00110001011001";
		Trees_din <= x"00093a0c";
		wait for Clk_period;
		Addr <=  "00110001011010";
		Trees_din <= x"1400fd04";
		wait for Clk_period;
		Addr <=  "00110001011011";
		Trees_din <= x"002931b9";
		wait for Clk_period;
		Addr <=  "00110001011100";
		Trees_din <= x"1600c704";
		wait for Clk_period;
		Addr <=  "00110001011101";
		Trees_din <= x"fff231b9";
		wait for Clk_period;
		Addr <=  "00110001011110";
		Trees_din <= x"ff7d31b9";
		wait for Clk_period;
		Addr <=  "00110001011111";
		Trees_din <= x"1900a810";
		wait for Clk_period;
		Addr <=  "00110001100000";
		Trees_din <= x"19009208";
		wait for Clk_period;
		Addr <=  "00110001100001";
		Trees_din <= x"09005204";
		wait for Clk_period;
		Addr <=  "00110001100010";
		Trees_din <= x"004431b9";
		wait for Clk_period;
		Addr <=  "00110001100011";
		Trees_din <= x"000131b9";
		wait for Clk_period;
		Addr <=  "00110001100100";
		Trees_din <= x"0f001404";
		wait for Clk_period;
		Addr <=  "00110001100101";
		Trees_din <= x"ff9631b9";
		wait for Clk_period;
		Addr <=  "00110001100110";
		Trees_din <= x"fffd31b9";
		wait for Clk_period;
		Addr <=  "00110001100111";
		Trees_din <= x"00115708";
		wait for Clk_period;
		Addr <=  "00110001101000";
		Trees_din <= x"1f000004";
		wait for Clk_period;
		Addr <=  "00110001101001";
		Trees_din <= x"007431b9";
		wait for Clk_period;
		Addr <=  "00110001101010";
		Trees_din <= x"ffd031b9";
		wait for Clk_period;
		Addr <=  "00110001101011";
		Trees_din <= x"00161e04";
		wait for Clk_period;
		Addr <=  "00110001101100";
		Trees_din <= x"ffa231b9";
		wait for Clk_period;
		Addr <=  "00110001101101";
		Trees_din <= x"003731b9";
		wait for Clk_period;
		Addr <=  "00110001101110";
		Trees_din <= x"0105aa48";
		wait for Clk_period;
		Addr <=  "00110001101111";
		Trees_din <= x"1200f718";
		wait for Clk_period;
		Addr <=  "00110001110000";
		Trees_din <= x"06fc3d14";
		wait for Clk_period;
		Addr <=  "00110001110001";
		Trees_din <= x"0efdd208";
		wait for Clk_period;
		Addr <=  "00110001110010";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00110001110011";
		Trees_din <= x"005832fd";
		wait for Clk_period;
		Addr <=  "00110001110100";
		Trees_din <= x"ffd632fd";
		wait for Clk_period;
		Addr <=  "00110001110101";
		Trees_din <= x"1a009c04";
		wait for Clk_period;
		Addr <=  "00110001110110";
		Trees_din <= x"fffc32fd";
		wait for Clk_period;
		Addr <=  "00110001110111";
		Trees_din <= x"1900aa04";
		wait for Clk_period;
		Addr <=  "00110001111000";
		Trees_din <= x"ff7932fd";
		wait for Clk_period;
		Addr <=  "00110001111001";
		Trees_din <= x"ffdc32fd";
		wait for Clk_period;
		Addr <=  "00110001111010";
		Trees_din <= x"003132fd";
		wait for Clk_period;
		Addr <=  "00110001111011";
		Trees_din <= x"0d02b01c";
		wait for Clk_period;
		Addr <=  "00110001111100";
		Trees_din <= x"11028610";
		wait for Clk_period;
		Addr <=  "00110001111101";
		Trees_din <= x"09005408";
		wait for Clk_period;
		Addr <=  "00110001111110";
		Trees_din <= x"0f03a304";
		wait for Clk_period;
		Addr <=  "00110001111111";
		Trees_din <= x"fff632fd";
		wait for Clk_period;
		Addr <=  "00110010000000";
		Trees_din <= x"006a32fd";
		wait for Clk_period;
		Addr <=  "00110010000001";
		Trees_din <= x"1a00b404";
		wait for Clk_period;
		Addr <=  "00110010000010";
		Trees_din <= x"000632fd";
		wait for Clk_period;
		Addr <=  "00110010000011";
		Trees_din <= x"ffae32fd";
		wait for Clk_period;
		Addr <=  "00110010000100";
		Trees_din <= x"13014804";
		wait for Clk_period;
		Addr <=  "00110010000101";
		Trees_din <= x"ff8432fd";
		wait for Clk_period;
		Addr <=  "00110010000110";
		Trees_din <= x"10fab204";
		wait for Clk_period;
		Addr <=  "00110010000111";
		Trees_din <= x"002832fd";
		wait for Clk_period;
		Addr <=  "00110010001000";
		Trees_din <= x"ffe032fd";
		wait for Clk_period;
		Addr <=  "00110010001001";
		Trees_din <= x"0d03370c";
		wait for Clk_period;
		Addr <=  "00110010001010";
		Trees_din <= x"17001d04";
		wait for Clk_period;
		Addr <=  "00110010001011";
		Trees_din <= x"ffdc32fd";
		wait for Clk_period;
		Addr <=  "00110010001100";
		Trees_din <= x"00082f04";
		wait for Clk_period;
		Addr <=  "00110010001101";
		Trees_din <= x"008a32fd";
		wait for Clk_period;
		Addr <=  "00110010001110";
		Trees_din <= x"002532fd";
		wait for Clk_period;
		Addr <=  "00110010001111";
		Trees_din <= x"1601b304";
		wait for Clk_period;
		Addr <=  "00110010010000";
		Trees_din <= x"002232fd";
		wait for Clk_period;
		Addr <=  "00110010010001";
		Trees_din <= x"ff9c32fd";
		wait for Clk_period;
		Addr <=  "00110010010010";
		Trees_din <= x"0d00051c";
		wait for Clk_period;
		Addr <=  "00110010010011";
		Trees_din <= x"1a00b810";
		wait for Clk_period;
		Addr <=  "00110010010100";
		Trees_din <= x"10027404";
		wait for Clk_period;
		Addr <=  "00110010010101";
		Trees_din <= x"ffac32fd";
		wait for Clk_period;
		Addr <=  "00110010010110";
		Trees_din <= x"1d005108";
		wait for Clk_period;
		Addr <=  "00110010010111";
		Trees_din <= x"0ef99404";
		wait for Clk_period;
		Addr <=  "00110010011000";
		Trees_din <= x"002032fd";
		wait for Clk_period;
		Addr <=  "00110010011001";
		Trees_din <= x"008032fd";
		wait for Clk_period;
		Addr <=  "00110010011010";
		Trees_din <= x"ffea32fd";
		wait for Clk_period;
		Addr <=  "00110010011011";
		Trees_din <= x"11028708";
		wait for Clk_period;
		Addr <=  "00110010011100";
		Trees_din <= x"0c00ed04";
		wait for Clk_period;
		Addr <=  "00110010011101";
		Trees_din <= x"ff7732fd";
		wait for Clk_period;
		Addr <=  "00110010011110";
		Trees_din <= x"ffe232fd";
		wait for Clk_period;
		Addr <=  "00110010011111";
		Trees_din <= x"fff832fd";
		wait for Clk_period;
		Addr <=  "00110010100000";
		Trees_din <= x"05fbaf20";
		wait for Clk_period;
		Addr <=  "00110010100001";
		Trees_din <= x"05fb6b10";
		wait for Clk_period;
		Addr <=  "00110010100010";
		Trees_din <= x"09005808";
		wait for Clk_period;
		Addr <=  "00110010100011";
		Trees_din <= x"11032704";
		wait for Clk_period;
		Addr <=  "00110010100100";
		Trees_din <= x"001632fd";
		wait for Clk_period;
		Addr <=  "00110010100101";
		Trees_din <= x"ffe432fd";
		wait for Clk_period;
		Addr <=  "00110010100110";
		Trees_din <= x"1102c004";
		wait for Clk_period;
		Addr <=  "00110010100111";
		Trees_din <= x"ffc432fd";
		wait for Clk_period;
		Addr <=  "00110010101000";
		Trees_din <= x"004232fd";
		wait for Clk_period;
		Addr <=  "00110010101001";
		Trees_din <= x"010c4908";
		wait for Clk_period;
		Addr <=  "00110010101010";
		Trees_din <= x"03fde004";
		wait for Clk_period;
		Addr <=  "00110010101011";
		Trees_din <= x"ff7d32fd";
		wait for Clk_period;
		Addr <=  "00110010101100";
		Trees_din <= x"fff132fd";
		wait for Clk_period;
		Addr <=  "00110010101101";
		Trees_din <= x"0e025a04";
		wait for Clk_period;
		Addr <=  "00110010101110";
		Trees_din <= x"ffc032fd";
		wait for Clk_period;
		Addr <=  "00110010101111";
		Trees_din <= x"005532fd";
		wait for Clk_period;
		Addr <=  "00110010110000";
		Trees_din <= x"0d024910";
		wait for Clk_period;
		Addr <=  "00110010110001";
		Trees_din <= x"09005508";
		wait for Clk_period;
		Addr <=  "00110010110010";
		Trees_din <= x"1004ee04";
		wait for Clk_period;
		Addr <=  "00110010110011";
		Trees_din <= x"001c32fd";
		wait for Clk_period;
		Addr <=  "00110010110100";
		Trees_din <= x"ffb632fd";
		wait for Clk_period;
		Addr <=  "00110010110101";
		Trees_din <= x"0f002b04";
		wait for Clk_period;
		Addr <=  "00110010110110";
		Trees_din <= x"fff232fd";
		wait for Clk_period;
		Addr <=  "00110010110111";
		Trees_din <= x"007c32fd";
		wait for Clk_period;
		Addr <=  "00110010111000";
		Trees_din <= x"20040008";
		wait for Clk_period;
		Addr <=  "00110010111001";
		Trees_din <= x"19008e04";
		wait for Clk_period;
		Addr <=  "00110010111010";
		Trees_din <= x"001532fd";
		wait for Clk_period;
		Addr <=  "00110010111011";
		Trees_din <= x"ff8132fd";
		wait for Clk_period;
		Addr <=  "00110010111100";
		Trees_din <= x"15009004";
		wait for Clk_period;
		Addr <=  "00110010111101";
		Trees_din <= x"ffbc32fd";
		wait for Clk_period;
		Addr <=  "00110010111110";
		Trees_din <= x"002732fd";
		wait for Clk_period;
		Addr <=  "00110010111111";
		Trees_din <= x"010a1f40";
		wait for Clk_period;
		Addr <=  "00110011000000";
		Trees_din <= x"13014d28";
		wait for Clk_period;
		Addr <=  "00110011000001";
		Trees_din <= x"15009914";
		wait for Clk_period;
		Addr <=  "00110011000010";
		Trees_din <= x"18003e04";
		wait for Clk_period;
		Addr <=  "00110011000011";
		Trees_din <= x"00743419";
		wait for Clk_period;
		Addr <=  "00110011000100";
		Trees_din <= x"06f98d08";
		wait for Clk_period;
		Addr <=  "00110011000101";
		Trees_din <= x"0afa1a04";
		wait for Clk_period;
		Addr <=  "00110011000110";
		Trees_din <= x"003b3419";
		wait for Clk_period;
		Addr <=  "00110011000111";
		Trees_din <= x"ffe93419";
		wait for Clk_period;
		Addr <=  "00110011001000";
		Trees_din <= x"0103f604";
		wait for Clk_period;
		Addr <=  "00110011001001";
		Trees_din <= x"ffc93419";
		wait for Clk_period;
		Addr <=  "00110011001010";
		Trees_din <= x"006a3419";
		wait for Clk_period;
		Addr <=  "00110011001011";
		Trees_din <= x"11fdc204";
		wait for Clk_period;
		Addr <=  "00110011001100";
		Trees_din <= x"00553419";
		wait for Clk_period;
		Addr <=  "00110011001101";
		Trees_din <= x"11021508";
		wait for Clk_period;
		Addr <=  "00110011001110";
		Trees_din <= x"14001b04";
		wait for Clk_period;
		Addr <=  "00110011001111";
		Trees_din <= x"00453419";
		wait for Clk_period;
		Addr <=  "00110011010000";
		Trees_din <= x"ffaa3419";
		wait for Clk_period;
		Addr <=  "00110011010001";
		Trees_din <= x"17026e04";
		wait for Clk_period;
		Addr <=  "00110011010010";
		Trees_din <= x"ffe53419";
		wait for Clk_period;
		Addr <=  "00110011010011";
		Trees_din <= x"003f3419";
		wait for Clk_period;
		Addr <=  "00110011010100";
		Trees_din <= x"06f35808";
		wait for Clk_period;
		Addr <=  "00110011010101";
		Trees_din <= x"0f016e04";
		wait for Clk_period;
		Addr <=  "00110011010110";
		Trees_din <= x"ffe33419";
		wait for Clk_period;
		Addr <=  "00110011010111";
		Trees_din <= x"00523419";
		wait for Clk_period;
		Addr <=  "00110011011000";
		Trees_din <= x"1d004e08";
		wait for Clk_period;
		Addr <=  "00110011011001";
		Trees_din <= x"02ffa304";
		wait for Clk_period;
		Addr <=  "00110011011010";
		Trees_din <= x"ffdd3419";
		wait for Clk_period;
		Addr <=  "00110011011011";
		Trees_din <= x"ff793419";
		wait for Clk_period;
		Addr <=  "00110011011100";
		Trees_din <= x"1b004704";
		wait for Clk_period;
		Addr <=  "00110011011101";
		Trees_din <= x"003a3419";
		wait for Clk_period;
		Addr <=  "00110011011110";
		Trees_din <= x"ffc83419";
		wait for Clk_period;
		Addr <=  "00110011011111";
		Trees_din <= x"020b0138";
		wait for Clk_period;
		Addr <=  "00110011100000";
		Trees_din <= x"0007fa1c";
		wait for Clk_period;
		Addr <=  "00110011100001";
		Trees_din <= x"1900a110";
		wait for Clk_period;
		Addr <=  "00110011100010";
		Trees_din <= x"07005c08";
		wait for Clk_period;
		Addr <=  "00110011100011";
		Trees_din <= x"00fda604";
		wait for Clk_period;
		Addr <=  "00110011100100";
		Trees_din <= x"ffe53419";
		wait for Clk_period;
		Addr <=  "00110011100101";
		Trees_din <= x"006d3419";
		wait for Clk_period;
		Addr <=  "00110011100110";
		Trees_din <= x"1a00b104";
		wait for Clk_period;
		Addr <=  "00110011100111";
		Trees_din <= x"ffb03419";
		wait for Clk_period;
		Addr <=  "00110011101000";
		Trees_din <= x"00233419";
		wait for Clk_period;
		Addr <=  "00110011101001";
		Trees_din <= x"09005104";
		wait for Clk_period;
		Addr <=  "00110011101010";
		Trees_din <= x"00623419";
		wait for Clk_period;
		Addr <=  "00110011101011";
		Trees_din <= x"0202a004";
		wait for Clk_period;
		Addr <=  "00110011101100";
		Trees_din <= x"00193419";
		wait for Clk_period;
		Addr <=  "00110011101101";
		Trees_din <= x"ffa33419";
		wait for Clk_period;
		Addr <=  "00110011101110";
		Trees_din <= x"00093a0c";
		wait for Clk_period;
		Addr <=  "00110011101111";
		Trees_din <= x"1400fd04";
		wait for Clk_period;
		Addr <=  "00110011110000";
		Trees_din <= x"003a3419";
		wait for Clk_period;
		Addr <=  "00110011110001";
		Trees_din <= x"1600c704";
		wait for Clk_period;
		Addr <=  "00110011110010";
		Trees_din <= x"fff73419";
		wait for Clk_period;
		Addr <=  "00110011110011";
		Trees_din <= x"ff893419";
		wait for Clk_period;
		Addr <=  "00110011110100";
		Trees_din <= x"0802b408";
		wait for Clk_period;
		Addr <=  "00110011110101";
		Trees_din <= x"08026904";
		wait for Clk_period;
		Addr <=  "00110011110110";
		Trees_din <= x"00083419";
		wait for Clk_period;
		Addr <=  "00110011110111";
		Trees_din <= x"ffa23419";
		wait for Clk_period;
		Addr <=  "00110011111000";
		Trees_din <= x"06f3b404";
		wait for Clk_period;
		Addr <=  "00110011111001";
		Trees_din <= x"ffc83419";
		wait for Clk_period;
		Addr <=  "00110011111010";
		Trees_din <= x"00473419";
		wait for Clk_period;
		Addr <=  "00110011111011";
		Trees_din <= x"0c019508";
		wait for Clk_period;
		Addr <=  "00110011111100";
		Trees_din <= x"10fade04";
		wait for Clk_period;
		Addr <=  "00110011111101";
		Trees_din <= x"ffdf3419";
		wait for Clk_period;
		Addr <=  "00110011111110";
		Trees_din <= x"ff903419";
		wait for Clk_period;
		Addr <=  "00110011111111";
		Trees_din <= x"15009708";
		wait for Clk_period;
		Addr <=  "00110100000000";
		Trees_din <= x"18004a04";
		wait for Clk_period;
		Addr <=  "00110100000001";
		Trees_din <= x"ff9f3419";
		wait for Clk_period;
		Addr <=  "00110100000010";
		Trees_din <= x"001e3419";
		wait for Clk_period;
		Addr <=  "00110100000011";
		Trees_din <= x"16020f04";
		wait for Clk_period;
		Addr <=  "00110100000100";
		Trees_din <= x"00023419";
		wait for Clk_period;
		Addr <=  "00110100000101";
		Trees_din <= x"005d3419";
		wait for Clk_period;
		Addr <=  "00110100000110";
		Trees_din <= x"0113e93c";
		wait for Clk_period;
		Addr <=  "00110100000111";
		Trees_din <= x"12fc6f0c";
		wait for Clk_period;
		Addr <=  "00110100001000";
		Trees_din <= x"0400ad08";
		wait for Clk_period;
		Addr <=  "00110100001001";
		Trees_din <= x"10020304";
		wait for Clk_period;
		Addr <=  "00110100001010";
		Trees_din <= x"ffea34bd";
		wait for Clk_period;
		Addr <=  "00110100001011";
		Trees_din <= x"ff9434bd";
		wait for Clk_period;
		Addr <=  "00110100001100";
		Trees_din <= x"001b34bd";
		wait for Clk_period;
		Addr <=  "00110100001101";
		Trees_din <= x"12fdae14";
		wait for Clk_period;
		Addr <=  "00110100001110";
		Trees_din <= x"02000008";
		wait for Clk_period;
		Addr <=  "00110100001111";
		Trees_din <= x"1a00d104";
		wait for Clk_period;
		Addr <=  "00110100010000";
		Trees_din <= x"ffc434bd";
		wait for Clk_period;
		Addr <=  "00110100010001";
		Trees_din <= x"001234bd";
		wait for Clk_period;
		Addr <=  "00110100010010";
		Trees_din <= x"02015404";
		wait for Clk_period;
		Addr <=  "00110100010011";
		Trees_din <= x"006c34bd";
		wait for Clk_period;
		Addr <=  "00110100010100";
		Trees_din <= x"17009804";
		wait for Clk_period;
		Addr <=  "00110100010101";
		Trees_din <= x"003034bd";
		wait for Clk_period;
		Addr <=  "00110100010110";
		Trees_din <= x"ffc134bd";
		wait for Clk_period;
		Addr <=  "00110100010111";
		Trees_din <= x"12fe290c";
		wait for Clk_period;
		Addr <=  "00110100011000";
		Trees_din <= x"010a6b04";
		wait for Clk_period;
		Addr <=  "00110100011001";
		Trees_din <= x"ff8434bd";
		wait for Clk_period;
		Addr <=  "00110100011010";
		Trees_din <= x"0a019904";
		wait for Clk_period;
		Addr <=  "00110100011011";
		Trees_din <= x"004534bd";
		wait for Clk_period;
		Addr <=  "00110100011100";
		Trees_din <= x"ffb034bd";
		wait for Clk_period;
		Addr <=  "00110100011101";
		Trees_din <= x"1403c008";
		wait for Clk_period;
		Addr <=  "00110100011110";
		Trees_din <= x"0f038404";
		wait for Clk_period;
		Addr <=  "00110100011111";
		Trees_din <= x"000134bd";
		wait for Clk_period;
		Addr <=  "00110100100000";
		Trees_din <= x"ffcc34bd";
		wait for Clk_period;
		Addr <=  "00110100100001";
		Trees_din <= x"0d000e04";
		wait for Clk_period;
		Addr <=  "00110100100010";
		Trees_din <= x"ffe834bd";
		wait for Clk_period;
		Addr <=  "00110100100011";
		Trees_din <= x"003334bd";
		wait for Clk_period;
		Addr <=  "00110100100100";
		Trees_din <= x"1e005e08";
		wait for Clk_period;
		Addr <=  "00110100100101";
		Trees_din <= x"01159304";
		wait for Clk_period;
		Addr <=  "00110100100110";
		Trees_din <= x"ffc134bd";
		wait for Clk_period;
		Addr <=  "00110100100111";
		Trees_din <= x"001f34bd";
		wait for Clk_period;
		Addr <=  "00110100101000";
		Trees_din <= x"00148708";
		wait for Clk_period;
		Addr <=  "00110100101001";
		Trees_din <= x"19008204";
		wait for Clk_period;
		Addr <=  "00110100101010";
		Trees_din <= x"000f34bd";
		wait for Clk_period;
		Addr <=  "00110100101011";
		Trees_din <= x"007334bd";
		wait for Clk_period;
		Addr <=  "00110100101100";
		Trees_din <= x"14014604";
		wait for Clk_period;
		Addr <=  "00110100101101";
		Trees_din <= x"002334bd";
		wait for Clk_period;
		Addr <=  "00110100101110";
		Trees_din <= x"ffd434bd";
		wait for Clk_period;
		Addr <=  "00110100101111";
		Trees_din <= x"010db654";
		wait for Clk_period;
		Addr <=  "00110100110000";
		Trees_din <= x"1400c128";
		wait for Clk_period;
		Addr <=  "00110100110001";
		Trees_din <= x"11fee80c";
		wait for Clk_period;
		Addr <=  "00110100110010";
		Trees_din <= x"1a00da08";
		wait for Clk_period;
		Addr <=  "00110100110011";
		Trees_din <= x"0f005e04";
		wait for Clk_period;
		Addr <=  "00110100110100";
		Trees_din <= x"ffcd35e1";
		wait for Clk_period;
		Addr <=  "00110100110101";
		Trees_din <= x"003e35e1";
		wait for Clk_period;
		Addr <=  "00110100110110";
		Trees_din <= x"006535e1";
		wait for Clk_period;
		Addr <=  "00110100110111";
		Trees_din <= x"05fa7c10";
		wait for Clk_period;
		Addr <=  "00110100111000";
		Trees_din <= x"0f000308";
		wait for Clk_period;
		Addr <=  "00110100111001";
		Trees_din <= x"0800af04";
		wait for Clk_period;
		Addr <=  "00110100111010";
		Trees_din <= x"004c35e1";
		wait for Clk_period;
		Addr <=  "00110100111011";
		Trees_din <= x"ffe335e1";
		wait for Clk_period;
		Addr <=  "00110100111100";
		Trees_din <= x"01061e04";
		wait for Clk_period;
		Addr <=  "00110100111101";
		Trees_din <= x"000935e1";
		wait for Clk_period;
		Addr <=  "00110100111110";
		Trees_din <= x"ff7c35e1";
		wait for Clk_period;
		Addr <=  "00110100111111";
		Trees_din <= x"05faab04";
		wait for Clk_period;
		Addr <=  "00110101000000";
		Trees_din <= x"005835e1";
		wait for Clk_period;
		Addr <=  "00110101000001";
		Trees_din <= x"0afabc04";
		wait for Clk_period;
		Addr <=  "00110101000010";
		Trees_din <= x"002335e1";
		wait for Clk_period;
		Addr <=  "00110101000011";
		Trees_din <= x"ffc535e1";
		wait for Clk_period;
		Addr <=  "00110101000100";
		Trees_din <= x"1702c81c";
		wait for Clk_period;
		Addr <=  "00110101000101";
		Trees_din <= x"16036810";
		wait for Clk_period;
		Addr <=  "00110101000110";
		Trees_din <= x"14027c08";
		wait for Clk_period;
		Addr <=  "00110101000111";
		Trees_din <= x"07005a04";
		wait for Clk_period;
		Addr <=  "00110101001000";
		Trees_din <= x"001e35e1";
		wait for Clk_period;
		Addr <=  "00110101001001";
		Trees_din <= x"ffd535e1";
		wait for Clk_period;
		Addr <=  "00110101001010";
		Trees_din <= x"0d024904";
		wait for Clk_period;
		Addr <=  "00110101001011";
		Trees_din <= x"fffe35e1";
		wait for Clk_period;
		Addr <=  "00110101001100";
		Trees_din <= x"ff9f35e1";
		wait for Clk_period;
		Addr <=  "00110101001101";
		Trees_din <= x"05f97c04";
		wait for Clk_period;
		Addr <=  "00110101001110";
		Trees_din <= x"002f35e1";
		wait for Clk_period;
		Addr <=  "00110101001111";
		Trees_din <= x"08027004";
		wait for Clk_period;
		Addr <=  "00110101010000";
		Trees_din <= x"ff7b35e1";
		wait for Clk_period;
		Addr <=  "00110101010001";
		Trees_din <= x"ffe235e1";
		wait for Clk_period;
		Addr <=  "00110101010010";
		Trees_din <= x"08004204";
		wait for Clk_period;
		Addr <=  "00110101010011";
		Trees_din <= x"ffd535e1";
		wait for Clk_period;
		Addr <=  "00110101010100";
		Trees_din <= x"17036008";
		wait for Clk_period;
		Addr <=  "00110101010101";
		Trees_din <= x"07005704";
		wait for Clk_period;
		Addr <=  "00110101010110";
		Trees_din <= x"007c35e1";
		wait for Clk_period;
		Addr <=  "00110101010111";
		Trees_din <= x"000f35e1";
		wait for Clk_period;
		Addr <=  "00110101011000";
		Trees_din <= x"ffea35e1";
		wait for Clk_period;
		Addr <=  "00110101011001";
		Trees_din <= x"21000034";
		wait for Clk_period;
		Addr <=  "00110101011010";
		Trees_din <= x"0e015f1c";
		wait for Clk_period;
		Addr <=  "00110101011011";
		Trees_din <= x"1800390c";
		wait for Clk_period;
		Addr <=  "00110101011100";
		Trees_din <= x"0803ae08";
		wait for Clk_period;
		Addr <=  "00110101011101";
		Trees_din <= x"000bca04";
		wait for Clk_period;
		Addr <=  "00110101011110";
		Trees_din <= x"ffe335e1";
		wait for Clk_period;
		Addr <=  "00110101011111";
		Trees_din <= x"ff8e35e1";
		wait for Clk_period;
		Addr <=  "00110101100000";
		Trees_din <= x"002935e1";
		wait for Clk_period;
		Addr <=  "00110101100001";
		Trees_din <= x"1b004808";
		wait for Clk_period;
		Addr <=  "00110101100010";
		Trees_din <= x"0c01ec04";
		wait for Clk_period;
		Addr <=  "00110101100011";
		Trees_din <= x"003635e1";
		wait for Clk_period;
		Addr <=  "00110101100100";
		Trees_din <= x"ffee35e1";
		wait for Clk_period;
		Addr <=  "00110101100101";
		Trees_din <= x"1a009804";
		wait for Clk_period;
		Addr <=  "00110101100110";
		Trees_din <= x"000c35e1";
		wait for Clk_period;
		Addr <=  "00110101100111";
		Trees_din <= x"ffa135e1";
		wait for Clk_period;
		Addr <=  "00110101101000";
		Trees_din <= x"11013d08";
		wait for Clk_period;
		Addr <=  "00110101101001";
		Trees_din <= x"12005e04";
		wait for Clk_period;
		Addr <=  "00110101101010";
		Trees_din <= x"002435e1";
		wait for Clk_period;
		Addr <=  "00110101101011";
		Trees_din <= x"008435e1";
		wait for Clk_period;
		Addr <=  "00110101101100";
		Trees_din <= x"1500a408";
		wait for Clk_period;
		Addr <=  "00110101101101";
		Trees_din <= x"1a00ca04";
		wait for Clk_period;
		Addr <=  "00110101101110";
		Trees_din <= x"002635e1";
		wait for Clk_period;
		Addr <=  "00110101101111";
		Trees_din <= x"ffc435e1";
		wait for Clk_period;
		Addr <=  "00110101110000";
		Trees_din <= x"00135a04";
		wait for Clk_period;
		Addr <=  "00110101110001";
		Trees_din <= x"007735e1";
		wait for Clk_period;
		Addr <=  "00110101110010";
		Trees_din <= x"fff335e1";
		wait for Clk_period;
		Addr <=  "00110101110011";
		Trees_din <= x"0afb1304";
		wait for Clk_period;
		Addr <=  "00110101110100";
		Trees_din <= x"001835e1";
		wait for Clk_period;
		Addr <=  "00110101110101";
		Trees_din <= x"02050704";
		wait for Clk_period;
		Addr <=  "00110101110110";
		Trees_din <= x"ff9735e1";
		wait for Clk_period;
		Addr <=  "00110101110111";
		Trees_din <= x"fff235e1";
		wait for Clk_period;
		Addr <=  "00110101111000";
		Trees_din <= x"01164264";
		wait for Clk_period;
		Addr <=  "00110101111001";
		Trees_din <= x"00111734";
		wait for Clk_period;
		Addr <=  "00110101111010";
		Trees_din <= x"21000020";
		wait for Clk_period;
		Addr <=  "00110101111011";
		Trees_din <= x"05fcb210";
		wait for Clk_period;
		Addr <=  "00110101111100";
		Trees_din <= x"05fc5208";
		wait for Clk_period;
		Addr <=  "00110101111101";
		Trees_din <= x"01081404";
		wait for Clk_period;
		Addr <=  "00110101111110";
		Trees_din <= x"ffee36b5";
		wait for Clk_period;
		Addr <=  "00110101111111";
		Trees_din <= x"000f36b5";
		wait for Clk_period;
		Addr <=  "00110110000000";
		Trees_din <= x"0b028604";
		wait for Clk_period;
		Addr <=  "00110110000001";
		Trees_din <= x"000036b5";
		wait for Clk_period;
		Addr <=  "00110110000010";
		Trees_din <= x"006436b5";
		wait for Clk_period;
		Addr <=  "00110110000011";
		Trees_din <= x"12019d08";
		wait for Clk_period;
		Addr <=  "00110110000100";
		Trees_din <= x"12017404";
		wait for Clk_period;
		Addr <=  "00110110000101";
		Trees_din <= x"fff636b5";
		wait for Clk_period;
		Addr <=  "00110110000110";
		Trees_din <= x"006636b5";
		wait for Clk_period;
		Addr <=  "00110110000111";
		Trees_din <= x"010b5404";
		wait for Clk_period;
		Addr <=  "00110110001000";
		Trees_din <= x"ffa736b5";
		wait for Clk_period;
		Addr <=  "00110110001001";
		Trees_din <= x"003736b5";
		wait for Clk_period;
		Addr <=  "00110110001010";
		Trees_din <= x"04fea408";
		wait for Clk_period;
		Addr <=  "00110110001011";
		Trees_din <= x"05f84b04";
		wait for Clk_period;
		Addr <=  "00110110001100";
		Trees_din <= x"fffc36b5";
		wait for Clk_period;
		Addr <=  "00110110001101";
		Trees_din <= x"ff8e36b5";
		wait for Clk_period;
		Addr <=  "00110110001110";
		Trees_din <= x"01076004";
		wait for Clk_period;
		Addr <=  "00110110001111";
		Trees_din <= x"ffd236b5";
		wait for Clk_period;
		Addr <=  "00110110010000";
		Trees_din <= x"13ffaf04";
		wait for Clk_period;
		Addr <=  "00110110010001";
		Trees_din <= x"005e36b5";
		wait for Clk_period;
		Addr <=  "00110110010010";
		Trees_din <= x"ffdc36b5";
		wait for Clk_period;
		Addr <=  "00110110010011";
		Trees_din <= x"09005a20";
		wait for Clk_period;
		Addr <=  "00110110010100";
		Trees_din <= x"1a00c310";
		wait for Clk_period;
		Addr <=  "00110110010101";
		Trees_din <= x"010fd308";
		wait for Clk_period;
		Addr <=  "00110110010110";
		Trees_din <= x"09004f04";
		wait for Clk_period;
		Addr <=  "00110110010111";
		Trees_din <= x"fff636b5";
		wait for Clk_period;
		Addr <=  "00110110011000";
		Trees_din <= x"ff7636b5";
		wait for Clk_period;
		Addr <=  "00110110011001";
		Trees_din <= x"1e007a04";
		wait for Clk_period;
		Addr <=  "00110110011010";
		Trees_din <= x"002136b5";
		wait for Clk_period;
		Addr <=  "00110110011011";
		Trees_din <= x"ffaa36b5";
		wait for Clk_period;
		Addr <=  "00110110011100";
		Trees_din <= x"1e006c08";
		wait for Clk_period;
		Addr <=  "00110110011101";
		Trees_din <= x"19009804";
		wait for Clk_period;
		Addr <=  "00110110011110";
		Trees_din <= x"ffa136b5";
		wait for Clk_period;
		Addr <=  "00110110011111";
		Trees_din <= x"fffe36b5";
		wait for Clk_period;
		Addr <=  "00110110100000";
		Trees_din <= x"13ffde04";
		wait for Clk_period;
		Addr <=  "00110110100001";
		Trees_din <= x"001036b5";
		wait for Clk_period;
		Addr <=  "00110110100010";
		Trees_din <= x"006736b5";
		wait for Clk_period;
		Addr <=  "00110110100011";
		Trees_din <= x"06f52304";
		wait for Clk_period;
		Addr <=  "00110110100100";
		Trees_din <= x"ffe136b5";
		wait for Clk_period;
		Addr <=  "00110110100101";
		Trees_din <= x"07005a08";
		wait for Clk_period;
		Addr <=  "00110110100110";
		Trees_din <= x"06f69e04";
		wait for Clk_period;
		Addr <=  "00110110100111";
		Trees_din <= x"007336b5";
		wait for Clk_period;
		Addr <=  "00110110101000";
		Trees_din <= x"001836b5";
		wait for Clk_period;
		Addr <=  "00110110101001";
		Trees_din <= x"fff636b5";
		wait for Clk_period;
		Addr <=  "00110110101010";
		Trees_din <= x"06f36504";
		wait for Clk_period;
		Addr <=  "00110110101011";
		Trees_din <= x"000b36b5";
		wait for Clk_period;
		Addr <=  "00110110101100";
		Trees_din <= x"005136b5";
		wait for Clk_period;
		Addr <=  "00110110101101";
		Trees_din <= x"1f000064";
		wait for Clk_period;
		Addr <=  "00110110101110";
		Trees_din <= x"010d4f2c";
		wait for Clk_period;
		Addr <=  "00110110101111";
		Trees_din <= x"0010b118";
		wait for Clk_period;
		Addr <=  "00110110110000";
		Trees_din <= x"03f7b30c";
		wait for Clk_period;
		Addr <=  "00110110110001";
		Trees_din <= x"10fbbf04";
		wait for Clk_period;
		Addr <=  "00110110110010";
		Trees_din <= x"002537c1";
		wait for Clk_period;
		Addr <=  "00110110110011";
		Trees_din <= x"15008e04";
		wait for Clk_period;
		Addr <=  "00110110110100";
		Trees_din <= x"ffeb37c1";
		wait for Clk_period;
		Addr <=  "00110110110101";
		Trees_din <= x"ff9037c1";
		wait for Clk_period;
		Addr <=  "00110110110110";
		Trees_din <= x"010d2808";
		wait for Clk_period;
		Addr <=  "00110110110111";
		Trees_din <= x"1d004404";
		wait for Clk_period;
		Addr <=  "00110110111000";
		Trees_din <= x"fff937c1";
		wait for Clk_period;
		Addr <=  "00110110111001";
		Trees_din <= x"001737c1";
		wait for Clk_period;
		Addr <=  "00110110111010";
		Trees_din <= x"ffab37c1";
		wait for Clk_period;
		Addr <=  "00110110111011";
		Trees_din <= x"1800430c";
		wait for Clk_period;
		Addr <=  "00110110111100";
		Trees_din <= x"1900a208";
		wait for Clk_period;
		Addr <=  "00110110111101";
		Trees_din <= x"1d004204";
		wait for Clk_period;
		Addr <=  "00110110111110";
		Trees_din <= x"003e37c1";
		wait for Clk_period;
		Addr <=  "00110110111111";
		Trees_din <= x"ffd737c1";
		wait for Clk_period;
		Addr <=  "00110111000000";
		Trees_din <= x"ffac37c1";
		wait for Clk_period;
		Addr <=  "00110111000001";
		Trees_din <= x"1c003704";
		wait for Clk_period;
		Addr <=  "00110111000010";
		Trees_din <= x"ffea37c1";
		wait for Clk_period;
		Addr <=  "00110111000011";
		Trees_din <= x"ff8337c1";
		wait for Clk_period;
		Addr <=  "00110111000100";
		Trees_din <= x"13001320";
		wait for Clk_period;
		Addr <=  "00110111000101";
		Trees_din <= x"0a028810";
		wait for Clk_period;
		Addr <=  "00110111000110";
		Trees_din <= x"0200d808";
		wait for Clk_period;
		Addr <=  "00110111000111";
		Trees_din <= x"00119204";
		wait for Clk_period;
		Addr <=  "00110111001000";
		Trees_din <= x"006337c1";
		wait for Clk_period;
		Addr <=  "00110111001001";
		Trees_din <= x"ffee37c1";
		wait for Clk_period;
		Addr <=  "00110111001010";
		Trees_din <= x"02019d04";
		wait for Clk_period;
		Addr <=  "00110111001011";
		Trees_din <= x"ffc137c1";
		wait for Clk_period;
		Addr <=  "00110111001100";
		Trees_din <= x"001037c1";
		wait for Clk_period;
		Addr <=  "00110111001101";
		Trees_din <= x"00119208";
		wait for Clk_period;
		Addr <=  "00110111001110";
		Trees_din <= x"1c004004";
		wait for Clk_period;
		Addr <=  "00110111001111";
		Trees_din <= x"ffb437c1";
		wait for Clk_period;
		Addr <=  "00110111010000";
		Trees_din <= x"002837c1";
		wait for Clk_period;
		Addr <=  "00110111010001";
		Trees_din <= x"0204c204";
		wait for Clk_period;
		Addr <=  "00110111010010";
		Trees_din <= x"ffeb37c1";
		wait for Clk_period;
		Addr <=  "00110111010011";
		Trees_din <= x"004d37c1";
		wait for Clk_period;
		Addr <=  "00110111010100";
		Trees_din <= x"010fff0c";
		wait for Clk_period;
		Addr <=  "00110111010101";
		Trees_din <= x"06f7fc08";
		wait for Clk_period;
		Addr <=  "00110111010110";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00110111010111";
		Trees_din <= x"001e37c1";
		wait for Clk_period;
		Addr <=  "00110111011000";
		Trees_din <= x"007737c1";
		wait for Clk_period;
		Addr <=  "00110111011001";
		Trees_din <= x"ffec37c1";
		wait for Clk_period;
		Addr <=  "00110111011010";
		Trees_din <= x"00138a08";
		wait for Clk_period;
		Addr <=  "00110111011011";
		Trees_din <= x"01117e04";
		wait for Clk_period;
		Addr <=  "00110111011100";
		Trees_din <= x"ffe337c1";
		wait for Clk_period;
		Addr <=  "00110111011101";
		Trees_din <= x"006537c1";
		wait for Clk_period;
		Addr <=  "00110111011110";
		Trees_din <= x"ffb337c1";
		wait for Clk_period;
		Addr <=  "00110111011111";
		Trees_din <= x"06f6f114";
		wait for Clk_period;
		Addr <=  "00110111100000";
		Trees_din <= x"0b04ee10";
		wait for Clk_period;
		Addr <=  "00110111100001";
		Trees_din <= x"0700580c";
		wait for Clk_period;
		Addr <=  "00110111100010";
		Trees_din <= x"1b002804";
		wait for Clk_period;
		Addr <=  "00110111100011";
		Trees_din <= x"fffd37c1";
		wait for Clk_period;
		Addr <=  "00110111100100";
		Trees_din <= x"22000004";
		wait for Clk_period;
		Addr <=  "00110111100101";
		Trees_din <= x"ff7d37c1";
		wait for Clk_period;
		Addr <=  "00110111100110";
		Trees_din <= x"fff137c1";
		wait for Clk_period;
		Addr <=  "00110111100111";
		Trees_din <= x"001637c1";
		wait for Clk_period;
		Addr <=  "00110111101000";
		Trees_din <= x"002837c1";
		wait for Clk_period;
		Addr <=  "00110111101001";
		Trees_din <= x"0f006a08";
		wait for Clk_period;
		Addr <=  "00110111101010";
		Trees_din <= x"00090504";
		wait for Clk_period;
		Addr <=  "00110111101011";
		Trees_din <= x"004237c1";
		wait for Clk_period;
		Addr <=  "00110111101100";
		Trees_din <= x"ffa937c1";
		wait for Clk_period;
		Addr <=  "00110111101101";
		Trees_din <= x"01099e04";
		wait for Clk_period;
		Addr <=  "00110111101110";
		Trees_din <= x"000537c1";
		wait for Clk_period;
		Addr <=  "00110111101111";
		Trees_din <= x"006f37c1";
		wait for Clk_period;
		Addr <=  "00110111110000";
		Trees_din <= x"010a1f6c";
		wait for Clk_period;
		Addr <=  "00110111110001";
		Trees_din <= x"07005738";
		wait for Clk_period;
		Addr <=  "00110111110010";
		Trees_din <= x"03fde01c";
		wait for Clk_period;
		Addr <=  "00110111110011";
		Trees_din <= x"1600630c";
		wait for Clk_period;
		Addr <=  "00110111110100";
		Trees_din <= x"11027704";
		wait for Clk_period;
		Addr <=  "00110111110101";
		Trees_din <= x"ffc838fd";
		wait for Clk_period;
		Addr <=  "00110111110110";
		Trees_din <= x"12027804";
		wait for Clk_period;
		Addr <=  "00110111110111";
		Trees_din <= x"006238fd";
		wait for Clk_period;
		Addr <=  "00110111111000";
		Trees_din <= x"001738fd";
		wait for Clk_period;
		Addr <=  "00110111111001";
		Trees_din <= x"06f2e408";
		wait for Clk_period;
		Addr <=  "00110111111010";
		Trees_din <= x"1102a504";
		wait for Clk_period;
		Addr <=  "00110111111011";
		Trees_din <= x"ffcb38fd";
		wait for Clk_period;
		Addr <=  "00110111111100";
		Trees_din <= x"005038fd";
		wait for Clk_period;
		Addr <=  "00110111111101";
		Trees_din <= x"01096904";
		wait for Clk_period;
		Addr <=  "00110111111110";
		Trees_din <= x"ff7f38fd";
		wait for Clk_period;
		Addr <=  "00110111111111";
		Trees_din <= x"fffe38fd";
		wait for Clk_period;
		Addr <=  "00111000000000";
		Trees_din <= x"06f6cc10";
		wait for Clk_period;
		Addr <=  "00111000000001";
		Trees_din <= x"07004d08";
		wait for Clk_period;
		Addr <=  "00111000000010";
		Trees_din <= x"05fc6304";
		wait for Clk_period;
		Addr <=  "00111000000011";
		Trees_din <= x"ffe938fd";
		wait for Clk_period;
		Addr <=  "00111000000100";
		Trees_din <= x"005338fd";
		wait for Clk_period;
		Addr <=  "00111000000101";
		Trees_din <= x"0d032204";
		wait for Clk_period;
		Addr <=  "00111000000110";
		Trees_din <= x"ff9d38fd";
		wait for Clk_period;
		Addr <=  "00111000000111";
		Trees_din <= x"001c38fd";
		wait for Clk_period;
		Addr <=  "00111000001000";
		Trees_din <= x"12ff9804";
		wait for Clk_period;
		Addr <=  "00111000001001";
		Trees_din <= x"ffc438fd";
		wait for Clk_period;
		Addr <=  "00111000001010";
		Trees_din <= x"01079604";
		wait for Clk_period;
		Addr <=  "00111000001011";
		Trees_din <= x"005238fd";
		wait for Clk_period;
		Addr <=  "00111000001100";
		Trees_din <= x"ffd838fd";
		wait for Clk_period;
		Addr <=  "00111000001101";
		Trees_din <= x"07005714";
		wait for Clk_period;
		Addr <=  "00111000001110";
		Trees_din <= x"02017b08";
		wait for Clk_period;
		Addr <=  "00111000001111";
		Trees_din <= x"06f5d004";
		wait for Clk_period;
		Addr <=  "00111000010000";
		Trees_din <= x"001b38fd";
		wait for Clk_period;
		Addr <=  "00111000010001";
		Trees_din <= x"ffb438fd";
		wait for Clk_period;
		Addr <=  "00111000010010";
		Trees_din <= x"0e01b208";
		wait for Clk_period;
		Addr <=  "00111000010011";
		Trees_din <= x"08017904";
		wait for Clk_period;
		Addr <=  "00111000010100";
		Trees_din <= x"009238fd";
		wait for Clk_period;
		Addr <=  "00111000010101";
		Trees_din <= x"002238fd";
		wait for Clk_period;
		Addr <=  "00111000010110";
		Trees_din <= x"fff738fd";
		wait for Clk_period;
		Addr <=  "00111000010111";
		Trees_din <= x"12017410";
		wait for Clk_period;
		Addr <=  "00111000011000";
		Trees_din <= x"13fda308";
		wait for Clk_period;
		Addr <=  "00111000011001";
		Trees_din <= x"0401a504";
		wait for Clk_period;
		Addr <=  "00111000011010";
		Trees_din <= x"002938fd";
		wait for Clk_period;
		Addr <=  "00111000011011";
		Trees_din <= x"ffa338fd";
		wait for Clk_period;
		Addr <=  "00111000011100";
		Trees_din <= x"03024704";
		wait for Clk_period;
		Addr <=  "00111000011101";
		Trees_din <= x"ff9038fd";
		wait for Clk_period;
		Addr <=  "00111000011110";
		Trees_din <= x"fff838fd";
		wait for Clk_period;
		Addr <=  "00111000011111";
		Trees_din <= x"12039108";
		wait for Clk_period;
		Addr <=  "00111000100000";
		Trees_din <= x"1102fb04";
		wait for Clk_period;
		Addr <=  "00111000100001";
		Trees_din <= x"000538fd";
		wait for Clk_period;
		Addr <=  "00111000100010";
		Trees_din <= x"005e38fd";
		wait for Clk_period;
		Addr <=  "00111000100011";
		Trees_din <= x"0c034b04";
		wait for Clk_period;
		Addr <=  "00111000100100";
		Trees_din <= x"ff9d38fd";
		wait for Clk_period;
		Addr <=  "00111000100101";
		Trees_din <= x"000038fd";
		wait for Clk_period;
		Addr <=  "00111000100110";
		Trees_din <= x"020b0124";
		wait for Clk_period;
		Addr <=  "00111000100111";
		Trees_din <= x"0f000010";
		wait for Clk_period;
		Addr <=  "00111000101000";
		Trees_din <= x"19009708";
		wait for Clk_period;
		Addr <=  "00111000101001";
		Trees_din <= x"03f91104";
		wait for Clk_period;
		Addr <=  "00111000101010";
		Trees_din <= x"fff738fd";
		wait for Clk_period;
		Addr <=  "00111000101011";
		Trees_din <= x"004638fd";
		wait for Clk_period;
		Addr <=  "00111000101100";
		Trees_din <= x"07005704";
		wait for Clk_period;
		Addr <=  "00111000101101";
		Trees_din <= x"ffe838fd";
		wait for Clk_period;
		Addr <=  "00111000101110";
		Trees_din <= x"ff8638fd";
		wait for Clk_period;
		Addr <=  "00111000101111";
		Trees_din <= x"14001304";
		wait for Clk_period;
		Addr <=  "00111000110000";
		Trees_din <= x"ffa138fd";
		wait for Clk_period;
		Addr <=  "00111000110001";
		Trees_din <= x"05fa2d08";
		wait for Clk_period;
		Addr <=  "00111000110010";
		Trees_din <= x"09005804";
		wait for Clk_period;
		Addr <=  "00111000110011";
		Trees_din <= x"000d38fd";
		wait for Clk_period;
		Addr <=  "00111000110100";
		Trees_din <= x"ffcd38fd";
		wait for Clk_period;
		Addr <=  "00111000110101";
		Trees_din <= x"1700f604";
		wait for Clk_period;
		Addr <=  "00111000110110";
		Trees_din <= x"000e38fd";
		wait for Clk_period;
		Addr <=  "00111000110111";
		Trees_din <= x"004138fd";
		wait for Clk_period;
		Addr <=  "00111000111000";
		Trees_din <= x"0110bb0c";
		wait for Clk_period;
		Addr <=  "00111000111001";
		Trees_din <= x"020db704";
		wait for Clk_period;
		Addr <=  "00111000111010";
		Trees_din <= x"ff9a38fd";
		wait for Clk_period;
		Addr <=  "00111000111011";
		Trees_din <= x"15009804";
		wait for Clk_period;
		Addr <=  "00111000111100";
		Trees_din <= x"ffcc38fd";
		wait for Clk_period;
		Addr <=  "00111000111101";
		Trees_din <= x"002d38fd";
		wait for Clk_period;
		Addr <=  "00111000111110";
		Trees_din <= x"002138fd";
		wait for Clk_period;
		Addr <=  "00111000111111";
		Trees_din <= x"0105aa30";
		wait for Clk_period;
		Addr <=  "00111001000000";
		Trees_din <= x"1200f710";
		wait for Clk_period;
		Addr <=  "00111001000001";
		Trees_din <= x"06fc3d0c";
		wait for Clk_period;
		Addr <=  "00111001000010";
		Trees_din <= x"0efdd204";
		wait for Clk_period;
		Addr <=  "00111001000011";
		Trees_din <= x"00143a01";
		wait for Clk_period;
		Addr <=  "00111001000100";
		Trees_din <= x"1d004f04";
		wait for Clk_period;
		Addr <=  "00111001000101";
		Trees_din <= x"ff893a01";
		wait for Clk_period;
		Addr <=  "00111001000110";
		Trees_din <= x"fff13a01";
		wait for Clk_period;
		Addr <=  "00111001000111";
		Trees_din <= x"002a3a01";
		wait for Clk_period;
		Addr <=  "00111001001000";
		Trees_din <= x"1900910c";
		wait for Clk_period;
		Addr <=  "00111001001001";
		Trees_din <= x"12019d04";
		wait for Clk_period;
		Addr <=  "00111001001010";
		Trees_din <= x"00143a01";
		wait for Clk_period;
		Addr <=  "00111001001011";
		Trees_din <= x"13015e04";
		wait for Clk_period;
		Addr <=  "00111001001100";
		Trees_din <= x"ff973a01";
		wait for Clk_period;
		Addr <=  "00111001001101";
		Trees_din <= x"ffec3a01";
		wait for Clk_period;
		Addr <=  "00111001001110";
		Trees_din <= x"1d00450c";
		wait for Clk_period;
		Addr <=  "00111001001111";
		Trees_din <= x"1a00d704";
		wait for Clk_period;
		Addr <=  "00111001010000";
		Trees_din <= x"ff9f3a01";
		wait for Clk_period;
		Addr <=  "00111001010001";
		Trees_din <= x"1a00dd04";
		wait for Clk_period;
		Addr <=  "00111001010010";
		Trees_din <= x"00503a01";
		wait for Clk_period;
		Addr <=  "00111001010011";
		Trees_din <= x"ffe53a01";
		wait for Clk_period;
		Addr <=  "00111001010100";
		Trees_din <= x"11027804";
		wait for Clk_period;
		Addr <=  "00111001010101";
		Trees_din <= x"00743a01";
		wait for Clk_period;
		Addr <=  "00111001010110";
		Trees_din <= x"00083a01";
		wait for Clk_period;
		Addr <=  "00111001010111";
		Trees_din <= x"03000c30";
		wait for Clk_period;
		Addr <=  "00111001011000";
		Trees_din <= x"0d000514";
		wait for Clk_period;
		Addr <=  "00111001011001";
		Trees_din <= x"1a00b80c";
		wait for Clk_period;
		Addr <=  "00111001011010";
		Trees_din <= x"10027404";
		wait for Clk_period;
		Addr <=  "00111001011011";
		Trees_din <= x"ffb73a01";
		wait for Clk_period;
		Addr <=  "00111001011100";
		Trees_din <= x"09005904";
		wait for Clk_period;
		Addr <=  "00111001011101";
		Trees_din <= x"000a3a01";
		wait for Clk_period;
		Addr <=  "00111001011110";
		Trees_din <= x"00633a01";
		wait for Clk_period;
		Addr <=  "00111001011111";
		Trees_din <= x"010de904";
		wait for Clk_period;
		Addr <=  "00111001100000";
		Trees_din <= x"ff883a01";
		wait for Clk_period;
		Addr <=  "00111001100001";
		Trees_din <= x"ffe03a01";
		wait for Clk_period;
		Addr <=  "00111001100010";
		Trees_din <= x"0e052810";
		wait for Clk_period;
		Addr <=  "00111001100011";
		Trees_din <= x"03fd8408";
		wait for Clk_period;
		Addr <=  "00111001100100";
		Trees_din <= x"0bf95604";
		wait for Clk_period;
		Addr <=  "00111001100101";
		Trees_din <= x"ffd83a01";
		wait for Clk_period;
		Addr <=  "00111001100110";
		Trees_din <= x"00093a01";
		wait for Clk_period;
		Addr <=  "00111001100111";
		Trees_din <= x"14027c04";
		wait for Clk_period;
		Addr <=  "00111001101000";
		Trees_din <= x"000c3a01";
		wait for Clk_period;
		Addr <=  "00111001101001";
		Trees_din <= x"ff8b3a01";
		wait for Clk_period;
		Addr <=  "00111001101010";
		Trees_din <= x"01098504";
		wait for Clk_period;
		Addr <=  "00111001101011";
		Trees_din <= x"fff53a01";
		wait for Clk_period;
		Addr <=  "00111001101100";
		Trees_din <= x"13fe1b04";
		wait for Clk_period;
		Addr <=  "00111001101101";
		Trees_din <= x"00153a01";
		wait for Clk_period;
		Addr <=  "00111001101110";
		Trees_din <= x"00663a01";
		wait for Clk_period;
		Addr <=  "00111001101111";
		Trees_din <= x"0f007310";
		wait for Clk_period;
		Addr <=  "00111001110000";
		Trees_din <= x"1c003108";
		wait for Clk_period;
		Addr <=  "00111001110001";
		Trees_din <= x"0e009f04";
		wait for Clk_period;
		Addr <=  "00111001110010";
		Trees_din <= x"fff93a01";
		wait for Clk_period;
		Addr <=  "00111001110011";
		Trees_din <= x"ff963a01";
		wait for Clk_period;
		Addr <=  "00111001110100";
		Trees_din <= x"1c003804";
		wait for Clk_period;
		Addr <=  "00111001110101";
		Trees_din <= x"003e3a01";
		wait for Clk_period;
		Addr <=  "00111001110110";
		Trees_din <= x"fff53a01";
		wait for Clk_period;
		Addr <=  "00111001110111";
		Trees_din <= x"0e02b00c";
		wait for Clk_period;
		Addr <=  "00111001111000";
		Trees_din <= x"01064704";
		wait for Clk_period;
		Addr <=  "00111001111001";
		Trees_din <= x"fff83a01";
		wait for Clk_period;
		Addr <=  "00111001111010";
		Trees_din <= x"21000004";
		wait for Clk_period;
		Addr <=  "00111001111011";
		Trees_din <= x"005e3a01";
		wait for Clk_period;
		Addr <=  "00111001111100";
		Trees_din <= x"fffb3a01";
		wait for Clk_period;
		Addr <=  "00111001111101";
		Trees_din <= x"10fb1604";
		wait for Clk_period;
		Addr <=  "00111001111110";
		Trees_din <= x"ffcd3a01";
		wait for Clk_period;
		Addr <=  "00111001111111";
		Trees_din <= x"000e3a01";
		wait for Clk_period;
		Addr <=  "00111010000000";
		Trees_din <= x"01082a38";
		wait for Clk_period;
		Addr <=  "00111010000001";
		Trees_din <= x"07005d30";
		wait for Clk_period;
		Addr <=  "00111010000010";
		Trees_din <= x"0f03dc20";
		wait for Clk_period;
		Addr <=  "00111010000011";
		Trees_din <= x"0d02c810";
		wait for Clk_period;
		Addr <=  "00111010000100";
		Trees_din <= x"1a00e308";
		wait for Clk_period;
		Addr <=  "00111010000101";
		Trees_din <= x"17000004";
		wait for Clk_period;
		Addr <=  "00111010000110";
		Trees_din <= x"ffee3b3d";
		wait for Clk_period;
		Addr <=  "00111010000111";
		Trees_din <= x"ffa33b3d";
		wait for Clk_period;
		Addr <=  "00111010001000";
		Trees_din <= x"07005704";
		wait for Clk_period;
		Addr <=  "00111010001001";
		Trees_din <= x"ffe33b3d";
		wait for Clk_period;
		Addr <=  "00111010001010";
		Trees_din <= x"00453b3d";
		wait for Clk_period;
		Addr <=  "00111010001011";
		Trees_din <= x"0d032a08";
		wait for Clk_period;
		Addr <=  "00111010001100";
		Trees_din <= x"1c002f04";
		wait for Clk_period;
		Addr <=  "00111010001101";
		Trees_din <= x"ffd33b3d";
		wait for Clk_period;
		Addr <=  "00111010001110";
		Trees_din <= x"004e3b3d";
		wait for Clk_period;
		Addr <=  "00111010001111";
		Trees_din <= x"0009b104";
		wait for Clk_period;
		Addr <=  "00111010010000";
		Trees_din <= x"fffa3b3d";
		wait for Clk_period;
		Addr <=  "00111010010001";
		Trees_din <= x"ff8f3b3d";
		wait for Clk_period;
		Addr <=  "00111010010010";
		Trees_din <= x"0d001208";
		wait for Clk_period;
		Addr <=  "00111010010011";
		Trees_din <= x"04f94b04";
		wait for Clk_period;
		Addr <=  "00111010010100";
		Trees_din <= x"00353b3d";
		wait for Clk_period;
		Addr <=  "00111010010101";
		Trees_din <= x"ffa93b3d";
		wait for Clk_period;
		Addr <=  "00111010010110";
		Trees_din <= x"02028904";
		wait for Clk_period;
		Addr <=  "00111010010111";
		Trees_din <= x"00553b3d";
		wait for Clk_period;
		Addr <=  "00111010011000";
		Trees_din <= x"00073b3d";
		wait for Clk_period;
		Addr <=  "00111010011001";
		Trees_din <= x"01059504";
		wait for Clk_period;
		Addr <=  "00111010011010";
		Trees_din <= x"00173b3d";
		wait for Clk_period;
		Addr <=  "00111010011011";
		Trees_din <= x"00523b3d";
		wait for Clk_period;
		Addr <=  "00111010011100";
		Trees_din <= x"03fbf640";
		wait for Clk_period;
		Addr <=  "00111010011101";
		Trees_din <= x"06f64820";
		wait for Clk_period;
		Addr <=  "00111010011110";
		Trees_din <= x"1c003210";
		wait for Clk_period;
		Addr <=  "00111010011111";
		Trees_din <= x"0f009708";
		wait for Clk_period;
		Addr <=  "00111010100000";
		Trees_din <= x"1e005f04";
		wait for Clk_period;
		Addr <=  "00111010100001";
		Trees_din <= x"00313b3d";
		wait for Clk_period;
		Addr <=  "00111010100010";
		Trees_din <= x"ffc13b3d";
		wait for Clk_period;
		Addr <=  "00111010100011";
		Trees_din <= x"01123c04";
		wait for Clk_period;
		Addr <=  "00111010100100";
		Trees_din <= x"ffa03b3d";
		wait for Clk_period;
		Addr <=  "00111010100101";
		Trees_din <= x"00143b3d";
		wait for Clk_period;
		Addr <=  "00111010100110";
		Trees_din <= x"1b003508";
		wait for Clk_period;
		Addr <=  "00111010100111";
		Trees_din <= x"14013104";
		wait for Clk_period;
		Addr <=  "00111010101000";
		Trees_din <= x"00643b3d";
		wait for Clk_period;
		Addr <=  "00111010101001";
		Trees_din <= x"000f3b3d";
		wait for Clk_period;
		Addr <=  "00111010101010";
		Trees_din <= x"17000104";
		wait for Clk_period;
		Addr <=  "00111010101011";
		Trees_din <= x"001a3b3d";
		wait for Clk_period;
		Addr <=  "00111010101100";
		Trees_din <= x"ffe73b3d";
		wait for Clk_period;
		Addr <=  "00111010101101";
		Trees_din <= x"00100410";
		wait for Clk_period;
		Addr <=  "00111010101110";
		Trees_din <= x"0e03fb08";
		wait for Clk_period;
		Addr <=  "00111010101111";
		Trees_din <= x"0d000504";
		wait for Clk_period;
		Addr <=  "00111010110000";
		Trees_din <= x"ffcb3b3d";
		wait for Clk_period;
		Addr <=  "00111010110001";
		Trees_din <= x"004b3b3d";
		wait for Clk_period;
		Addr <=  "00111010110010";
		Trees_din <= x"14021e04";
		wait for Clk_period;
		Addr <=  "00111010110011";
		Trees_din <= x"ffad3b3d";
		wait for Clk_period;
		Addr <=  "00111010110100";
		Trees_din <= x"fff33b3d";
		wait for Clk_period;
		Addr <=  "00111010110101";
		Trees_din <= x"0e022208";
		wait for Clk_period;
		Addr <=  "00111010110110";
		Trees_din <= x"02062104";
		wait for Clk_period;
		Addr <=  "00111010110111";
		Trees_din <= x"ffbf3b3d";
		wait for Clk_period;
		Addr <=  "00111010111000";
		Trees_din <= x"00453b3d";
		wait for Clk_period;
		Addr <=  "00111010111001";
		Trees_din <= x"06f77e04";
		wait for Clk_period;
		Addr <=  "00111010111010";
		Trees_din <= x"005c3b3d";
		wait for Clk_period;
		Addr <=  "00111010111011";
		Trees_din <= x"ffe33b3d";
		wait for Clk_period;
		Addr <=  "00111010111100";
		Trees_din <= x"0900591c";
		wait for Clk_period;
		Addr <=  "00111010111101";
		Trees_din <= x"06f82e10";
		wait for Clk_period;
		Addr <=  "00111010111110";
		Trees_din <= x"0c00e308";
		wait for Clk_period;
		Addr <=  "00111010111111";
		Trees_din <= x"10028404";
		wait for Clk_period;
		Addr <=  "00111011000000";
		Trees_din <= x"ffbd3b3d";
		wait for Clk_period;
		Addr <=  "00111011000001";
		Trees_din <= x"00263b3d";
		wait for Clk_period;
		Addr <=  "00111011000010";
		Trees_din <= x"0b044d04";
		wait for Clk_period;
		Addr <=  "00111011000011";
		Trees_din <= x"00573b3d";
		wait for Clk_period;
		Addr <=  "00111011000100";
		Trees_din <= x"ffff3b3d";
		wait for Clk_period;
		Addr <=  "00111011000101";
		Trees_din <= x"05f88104";
		wait for Clk_period;
		Addr <=  "00111011000110";
		Trees_din <= x"00363b3d";
		wait for Clk_period;
		Addr <=  "00111011000111";
		Trees_din <= x"02016004";
		wait for Clk_period;
		Addr <=  "00111011001000";
		Trees_din <= x"00113b3d";
		wait for Clk_period;
		Addr <=  "00111011001001";
		Trees_din <= x"ff8b3b3d";
		wait for Clk_period;
		Addr <=  "00111011001010";
		Trees_din <= x"13ffe608";
		wait for Clk_period;
		Addr <=  "00111011001011";
		Trees_din <= x"13ff5804";
		wait for Clk_period;
		Addr <=  "00111011001100";
		Trees_din <= x"ff8f3b3d";
		wait for Clk_period;
		Addr <=  "00111011001101";
		Trees_din <= x"ffeb3b3d";
		wait for Clk_period;
		Addr <=  "00111011001110";
		Trees_din <= x"00463b3d";
		wait for Clk_period;
		Addr <=  "00111011001111";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  1
        -----------
		Addr <=  "00000000000000";
		Trees_din <= x"000e4f70";
		wait for Clk_period;
		Addr <=  "00000000000001";
		Trees_din <= x"00097434";
		wait for Clk_period;
		Addr <=  "00000000000010";
		Trees_din <= x"0003aa14";
		wait for Clk_period;
		Addr <=  "00000000000011";
		Trees_din <= x"1b006610";
		wait for Clk_period;
		Addr <=  "00000000000100";
		Trees_din <= x"1d005a08";
		wait for Clk_period;
		Addr <=  "00000000000101";
		Trees_din <= x"0000af04";
		wait for Clk_period;
		Addr <=  "00000000000110";
		Trees_din <= x"ff5601a5";
		wait for Clk_period;
		Addr <=  "00000000000111";
		Trees_din <= x"ff7701a5";
		wait for Clk_period;
		Addr <=  "00000000001000";
		Trees_din <= x"0d002a04";
		wait for Clk_period;
		Addr <=  "00000000001001";
		Trees_din <= x"013c01a5";
		wait for Clk_period;
		Addr <=  "00000000001010";
		Trees_din <= x"ff7001a5";
		wait for Clk_period;
		Addr <=  "00000000001011";
		Trees_din <= x"008e01a5";
		wait for Clk_period;
		Addr <=  "00000000001100";
		Trees_din <= x"03fe5110";
		wait for Clk_period;
		Addr <=  "00000000001101";
		Trees_din <= x"020b0108";
		wait for Clk_period;
		Addr <=  "00000000001110";
		Trees_din <= x"05fb0f04";
		wait for Clk_period;
		Addr <=  "00000000001111";
		Trees_din <= x"ff8b01a5";
		wait for Clk_period;
		Addr <=  "00000000010000";
		Trees_din <= x"003b01a5";
		wait for Clk_period;
		Addr <=  "00000000010001";
		Trees_din <= x"11047904";
		wait for Clk_period;
		Addr <=  "00000000010010";
		Trees_din <= x"ff5001a5";
		wait for Clk_period;
		Addr <=  "00000000010011";
		Trees_din <= x"ffd001a5";
		wait for Clk_period;
		Addr <=  "00000000010100";
		Trees_din <= x"0400f008";
		wait for Clk_period;
		Addr <=  "00000000010101";
		Trees_din <= x"06fa4504";
		wait for Clk_period;
		Addr <=  "00000000010110";
		Trees_din <= x"ffd101a5";
		wait for Clk_period;
		Addr <=  "00000000010111";
		Trees_din <= x"00d701a5";
		wait for Clk_period;
		Addr <=  "00000000011000";
		Trees_din <= x"05fe9604";
		wait for Clk_period;
		Addr <=  "00000000011001";
		Trees_din <= x"01d801a5";
		wait for Clk_period;
		Addr <=  "00000000011010";
		Trees_din <= x"ffd901a5";
		wait for Clk_period;
		Addr <=  "00000000011011";
		Trees_din <= x"03fa871c";
		wait for Clk_period;
		Addr <=  "00000000011100";
		Trees_din <= x"010ed010";
		wait for Clk_period;
		Addr <=  "00000000011101";
		Trees_din <= x"0208db08";
		wait for Clk_period;
		Addr <=  "00000000011110";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00000000011111";
		Trees_din <= x"020801a5";
		wait for Clk_period;
		Addr <=  "00000000100000";
		Trees_din <= x"007c01a5";
		wait for Clk_period;
		Addr <=  "00000000100001";
		Trees_din <= x"08000f04";
		wait for Clk_period;
		Addr <=  "00000000100010";
		Trees_din <= x"00c101a5";
		wait for Clk_period;
		Addr <=  "00000000100011";
		Trees_din <= x"ff9101a5";
		wait for Clk_period;
		Addr <=  "00000000100100";
		Trees_din <= x"01139008";
		wait for Clk_period;
		Addr <=  "00000000100101";
		Trees_din <= x"0afc8304";
		wait for Clk_period;
		Addr <=  "00000000100110";
		Trees_din <= x"ff7201a5";
		wait for Clk_period;
		Addr <=  "00000000100111";
		Trees_din <= x"004b01a5";
		wait for Clk_period;
		Addr <=  "00000000101000";
		Trees_din <= x"ff5601a5";
		wait for Clk_period;
		Addr <=  "00000000101001";
		Trees_din <= x"01090e10";
		wait for Clk_period;
		Addr <=  "00000000101010";
		Trees_din <= x"02068508";
		wait for Clk_period;
		Addr <=  "00000000101011";
		Trees_din <= x"07005c04";
		wait for Clk_period;
		Addr <=  "00000000101100";
		Trees_din <= x"038801a5";
		wait for Clk_period;
		Addr <=  "00000000101101";
		Trees_din <= x"00c101a5";
		wait for Clk_period;
		Addr <=  "00000000101110";
		Trees_din <= x"0103c204";
		wait for Clk_period;
		Addr <=  "00000000101111";
		Trees_din <= x"012001a5";
		wait for Clk_period;
		Addr <=  "00000000110000";
		Trees_din <= x"ffa701a5";
		wait for Clk_period;
		Addr <=  "00000000110001";
		Trees_din <= x"0afc8308";
		wait for Clk_period;
		Addr <=  "00000000110010";
		Trees_din <= x"0c004604";
		wait for Clk_period;
		Addr <=  "00000000110011";
		Trees_din <= x"002701a5";
		wait for Clk_period;
		Addr <=  "00000000110100";
		Trees_din <= x"ff6b01a5";
		wait for Clk_period;
		Addr <=  "00000000110101";
		Trees_din <= x"06f73004";
		wait for Clk_period;
		Addr <=  "00000000110110";
		Trees_din <= x"020201a5";
		wait for Clk_period;
		Addr <=  "00000000110111";
		Trees_din <= x"ff8101a5";
		wait for Clk_period;
		Addr <=  "00000000111000";
		Trees_din <= x"0111ec34";
		wait for Clk_period;
		Addr <=  "00000000111001";
		Trees_din <= x"0011ff20";
		wait for Clk_period;
		Addr <=  "00000000111010";
		Trees_din <= x"010aed10";
		wait for Clk_period;
		Addr <=  "00000000111011";
		Trees_din <= x"020abe08";
		wait for Clk_period;
		Addr <=  "00000000111100";
		Trees_din <= x"05f70004";
		wait for Clk_period;
		Addr <=  "00000000111101";
		Trees_din <= x"015401a5";
		wait for Clk_period;
		Addr <=  "00000000111110";
		Trees_din <= x"03c101a5";
		wait for Clk_period;
		Addr <=  "00000000111111";
		Trees_din <= x"0c026304";
		wait for Clk_period;
		Addr <=  "00000001000000";
		Trees_din <= x"017401a5";
		wait for Clk_period;
		Addr <=  "00000001000001";
		Trees_din <= x"000a01a5";
		wait for Clk_period;
		Addr <=  "00000001000010";
		Trees_din <= x"1500a308";
		wait for Clk_period;
		Addr <=  "00000001000011";
		Trees_din <= x"05fc8504";
		wait for Clk_period;
		Addr <=  "00000001000100";
		Trees_din <= x"026501a5";
		wait for Clk_period;
		Addr <=  "00000001000101";
		Trees_din <= x"ff9d01a5";
		wait for Clk_period;
		Addr <=  "00000001000110";
		Trees_din <= x"0f005504";
		wait for Clk_period;
		Addr <=  "00000001000111";
		Trees_din <= x"ffb001a5";
		wait for Clk_period;
		Addr <=  "00000001001000";
		Trees_din <= x"01c201a5";
		wait for Clk_period;
		Addr <=  "00000001001001";
		Trees_din <= x"00167610";
		wait for Clk_period;
		Addr <=  "00000001001010";
		Trees_din <= x"02097608";
		wait for Clk_period;
		Addr <=  "00000001001011";
		Trees_din <= x"0e052804";
		wait for Clk_period;
		Addr <=  "00000001001100";
		Trees_din <= x"03ea01a5";
		wait for Clk_period;
		Addr <=  "00000001001101";
		Trees_din <= x"019001a5";
		wait for Clk_period;
		Addr <=  "00000001001110";
		Trees_din <= x"09005904";
		wait for Clk_period;
		Addr <=  "00000001001111";
		Trees_din <= x"02dc01a5";
		wait for Clk_period;
		Addr <=  "00000001010000";
		Trees_din <= x"001601a5";
		wait for Clk_period;
		Addr <=  "00000001010001";
		Trees_din <= x"042f01a5";
		wait for Clk_period;
		Addr <=  "00000001010010";
		Trees_din <= x"0015001c";
		wait for Clk_period;
		Addr <=  "00000001010011";
		Trees_din <= x"0011ff0c";
		wait for Clk_period;
		Addr <=  "00000001010100";
		Trees_din <= x"0efa8a04";
		wait for Clk_period;
		Addr <=  "00000001010101";
		Trees_din <= x"01c601a5";
		wait for Clk_period;
		Addr <=  "00000001010110";
		Trees_din <= x"01139004";
		wait for Clk_period;
		Addr <=  "00000001010111";
		Trees_din <= x"001601a5";
		wait for Clk_period;
		Addr <=  "00000001011000";
		Trees_din <= x"ff5c01a5";
		wait for Clk_period;
		Addr <=  "00000001011001";
		Trees_din <= x"0114d608";
		wait for Clk_period;
		Addr <=  "00000001011010";
		Trees_din <= x"0c032b04";
		wait for Clk_period;
		Addr <=  "00000001011011";
		Trees_din <= x"021801a5";
		wait for Clk_period;
		Addr <=  "00000001011100";
		Trees_din <= x"002701a5";
		wait for Clk_period;
		Addr <=  "00000001011101";
		Trees_din <= x"02043f04";
		wait for Clk_period;
		Addr <=  "00000001011110";
		Trees_din <= x"00b201a5";
		wait for Clk_period;
		Addr <=  "00000001011111";
		Trees_din <= x"ff7d01a5";
		wait for Clk_period;
		Addr <=  "00000001100000";
		Trees_din <= x"0116420c";
		wait for Clk_period;
		Addr <=  "00000001100001";
		Trees_din <= x"00167608";
		wait for Clk_period;
		Addr <=  "00000001100010";
		Trees_din <= x"03f37e04";
		wait for Clk_period;
		Addr <=  "00000001100011";
		Trees_din <= x"005901a5";
		wait for Clk_period;
		Addr <=  "00000001100100";
		Trees_din <= x"028401a5";
		wait for Clk_period;
		Addr <=  "00000001100101";
		Trees_din <= x"03a701a5";
		wait for Clk_period;
		Addr <=  "00000001100110";
		Trees_din <= x"0b040404";
		wait for Clk_period;
		Addr <=  "00000001100111";
		Trees_din <= x"000001a5";
		wait for Clk_period;
		Addr <=  "00000001101000";
		Trees_din <= x"01c601a5";
		wait for Clk_period;
		Addr <=  "00000001101001";
		Trees_din <= x"000ceb60";
		wait for Clk_period;
		Addr <=  "00000001101010";
		Trees_din <= x"0004a124";
		wait for Clk_period;
		Addr <=  "00000001101011";
		Trees_din <= x"14000b08";
		wait for Clk_period;
		Addr <=  "00000001101100";
		Trees_din <= x"19008a04";
		wait for Clk_period;
		Addr <=  "00000001101101";
		Trees_din <= x"ff9802f1";
		wait for Clk_period;
		Addr <=  "00000001101110";
		Trees_din <= x"016e02f1";
		wait for Clk_period;
		Addr <=  "00000001101111";
		Trees_din <= x"0000af0c";
		wait for Clk_period;
		Addr <=  "00000001110000";
		Trees_din <= x"1204f608";
		wait for Clk_period;
		Addr <=  "00000001110001";
		Trees_din <= x"09003e04";
		wait for Clk_period;
		Addr <=  "00000001110010";
		Trees_din <= x"fff502f1";
		wait for Clk_period;
		Addr <=  "00000001110011";
		Trees_din <= x"ff5902f1";
		wait for Clk_period;
		Addr <=  "00000001110100";
		Trees_din <= x"002702f1";
		wait for Clk_period;
		Addr <=  "00000001110101";
		Trees_din <= x"03ff5408";
		wait for Clk_period;
		Addr <=  "00000001110110";
		Trees_din <= x"14001d04";
		wait for Clk_period;
		Addr <=  "00000001110111";
		Trees_din <= x"ffee02f1";
		wait for Clk_period;
		Addr <=  "00000001111000";
		Trees_din <= x"ff5402f1";
		wait for Clk_period;
		Addr <=  "00000001111001";
		Trees_din <= x"0402ab04";
		wait for Clk_period;
		Addr <=  "00000001111010";
		Trees_din <= x"ff7902f1";
		wait for Clk_period;
		Addr <=  "00000001111011";
		Trees_din <= x"004302f1";
		wait for Clk_period;
		Addr <=  "00000001111100";
		Trees_din <= x"03fa871c";
		wait for Clk_period;
		Addr <=  "00000001111101";
		Trees_din <= x"020abe10";
		wait for Clk_period;
		Addr <=  "00000001111110";
		Trees_din <= x"05fb0f08";
		wait for Clk_period;
		Addr <=  "00000001111111";
		Trees_din <= x"13019604";
		wait for Clk_period;
		Addr <=  "00000010000000";
		Trees_din <= x"ff7f02f1";
		wait for Clk_period;
		Addr <=  "00000010000001";
		Trees_din <= x"009c02f1";
		wait for Clk_period;
		Addr <=  "00000010000010";
		Trees_din <= x"09005004";
		wait for Clk_period;
		Addr <=  "00000010000011";
		Trees_din <= x"ff6802f1";
		wait for Clk_period;
		Addr <=  "00000010000100";
		Trees_din <= x"00da02f1";
		wait for Clk_period;
		Addr <=  "00000010000101";
		Trees_din <= x"06f6f104";
		wait for Clk_period;
		Addr <=  "00000010000110";
		Trees_din <= x"ff5702f1";
		wait for Clk_period;
		Addr <=  "00000010000111";
		Trees_din <= x"11007904";
		wait for Clk_period;
		Addr <=  "00000010001000";
		Trees_din <= x"00b602f1";
		wait for Clk_period;
		Addr <=  "00000010001001";
		Trees_din <= x"ff9802f1";
		wait for Clk_period;
		Addr <=  "00000010001010";
		Trees_din <= x"02077510";
		wait for Clk_period;
		Addr <=  "00000010001011";
		Trees_din <= x"010b5408";
		wait for Clk_period;
		Addr <=  "00000010001100";
		Trees_din <= x"05005804";
		wait for Clk_period;
		Addr <=  "00000010001101";
		Trees_din <= x"012902f1";
		wait for Clk_period;
		Addr <=  "00000010001110";
		Trees_din <= x"ffdb02f1";
		wait for Clk_period;
		Addr <=  "00000010001111";
		Trees_din <= x"03facd04";
		wait for Clk_period;
		Addr <=  "00000010010000";
		Trees_din <= x"015c02f1";
		wait for Clk_period;
		Addr <=  "00000010010001";
		Trees_din <= x"ffbe02f1";
		wait for Clk_period;
		Addr <=  "00000010010010";
		Trees_din <= x"0af7e808";
		wait for Clk_period;
		Addr <=  "00000010010011";
		Trees_din <= x"19008f04";
		wait for Clk_period;
		Addr <=  "00000010010100";
		Trees_din <= x"ff9f02f1";
		wait for Clk_period;
		Addr <=  "00000010010101";
		Trees_din <= x"018d02f1";
		wait for Clk_period;
		Addr <=  "00000010010110";
		Trees_din <= x"0b028004";
		wait for Clk_period;
		Addr <=  "00000010010111";
		Trees_din <= x"001e02f1";
		wait for Clk_period;
		Addr <=  "00000010011000";
		Trees_din <= x"ff5a02f1";
		wait for Clk_period;
		Addr <=  "00000010011001";
		Trees_din <= x"01159330";
		wait for Clk_period;
		Addr <=  "00000010011010";
		Trees_din <= x"000fd31c";
		wait for Clk_period;
		Addr <=  "00000010011011";
		Trees_din <= x"03f68f0c";
		wait for Clk_period;
		Addr <=  "00000010011100";
		Trees_din <= x"04fc5b08";
		wait for Clk_period;
		Addr <=  "00000010011101";
		Trees_din <= x"0d037f04";
		wait for Clk_period;
		Addr <=  "00000010011110";
		Trees_din <= x"ff7802f1";
		wait for Clk_period;
		Addr <=  "00000010011111";
		Trees_din <= x"007902f1";
		wait for Clk_period;
		Addr <=  "00000010100000";
		Trees_din <= x"010702f1";
		wait for Clk_period;
		Addr <=  "00000010100001";
		Trees_din <= x"01082a08";
		wait for Clk_period;
		Addr <=  "00000010100010";
		Trees_din <= x"0208db04";
		wait for Clk_period;
		Addr <=  "00000010100011";
		Trees_din <= x"01a102f1";
		wait for Clk_period;
		Addr <=  "00000010100100";
		Trees_din <= x"005902f1";
		wait for Clk_period;
		Addr <=  "00000010100101";
		Trees_din <= x"06f62e04";
		wait for Clk_period;
		Addr <=  "00000010100110";
		Trees_din <= x"013402f1";
		wait for Clk_period;
		Addr <=  "00000010100111";
		Trees_din <= x"005c02f1";
		wait for Clk_period;
		Addr <=  "00000010101000";
		Trees_din <= x"010d4f04";
		wait for Clk_period;
		Addr <=  "00000010101001";
		Trees_din <= x"01a802f1";
		wait for Clk_period;
		Addr <=  "00000010101010";
		Trees_din <= x"00135a08";
		wait for Clk_period;
		Addr <=  "00000010101011";
		Trees_din <= x"0c031c04";
		wait for Clk_period;
		Addr <=  "00000010101100";
		Trees_din <= x"013a02f1";
		wait for Clk_period;
		Addr <=  "00000010101101";
		Trees_din <= x"002d02f1";
		wait for Clk_period;
		Addr <=  "00000010101110";
		Trees_din <= x"0bf8e904";
		wait for Clk_period;
		Addr <=  "00000010101111";
		Trees_din <= x"004702f1";
		wait for Clk_period;
		Addr <=  "00000010110000";
		Trees_din <= x"019102f1";
		wait for Clk_period;
		Addr <=  "00000010110001";
		Trees_din <= x"0013bd04";
		wait for Clk_period;
		Addr <=  "00000010110010";
		Trees_din <= x"ff6202f1";
		wait for Clk_period;
		Addr <=  "00000010110011";
		Trees_din <= x"0afb1008";
		wait for Clk_period;
		Addr <=  "00000010110100";
		Trees_din <= x"07005a04";
		wait for Clk_period;
		Addr <=  "00000010110101";
		Trees_din <= x"ffa202f1";
		wait for Clk_period;
		Addr <=  "00000010110110";
		Trees_din <= x"002f02f1";
		wait for Clk_period;
		Addr <=  "00000010110111";
		Trees_din <= x"0b040408";
		wait for Clk_period;
		Addr <=  "00000010111000";
		Trees_din <= x"0d00e504";
		wait for Clk_period;
		Addr <=  "00000010111001";
		Trees_din <= x"013702f1";
		wait for Clk_period;
		Addr <=  "00000010111010";
		Trees_din <= x"ff9402f1";
		wait for Clk_period;
		Addr <=  "00000010111011";
		Trees_din <= x"01d502f1";
		wait for Clk_period;
		Addr <=  "00000010111100";
		Trees_din <= x"000bca70";
		wait for Clk_period;
		Addr <=  "00000010111101";
		Trees_din <= x"0004a134";
		wait for Clk_period;
		Addr <=  "00000010111110";
		Trees_din <= x"0000af14";
		wait for Clk_period;
		Addr <=  "00000010111111";
		Trees_din <= x"09003e08";
		wait for Clk_period;
		Addr <=  "00000011000000";
		Trees_din <= x"06f63b04";
		wait for Clk_period;
		Addr <=  "00000011000001";
		Trees_din <= x"ffa50485";
		wait for Clk_period;
		Addr <=  "00000011000010";
		Trees_din <= x"00c50485";
		wait for Clk_period;
		Addr <=  "00000011000011";
		Trees_din <= x"0803f908";
		wait for Clk_period;
		Addr <=  "00000011000100";
		Trees_din <= x"1204f604";
		wait for Clk_period;
		Addr <=  "00000011000101";
		Trees_din <= x"ff5e0485";
		wait for Clk_period;
		Addr <=  "00000011000110";
		Trees_din <= x"00290485";
		wait for Clk_period;
		Addr <=  "00000011000111";
		Trees_din <= x"002f0485";
		wait for Clk_period;
		Addr <=  "00000011001000";
		Trees_din <= x"04025d10";
		wait for Clk_period;
		Addr <=  "00000011001001";
		Trees_din <= x"0d03ae08";
		wait for Clk_period;
		Addr <=  "00000011001010";
		Trees_din <= x"0ef9a204";
		wait for Clk_period;
		Addr <=  "00000011001011";
		Trees_din <= x"ffc20485";
		wait for Clk_period;
		Addr <=  "00000011001100";
		Trees_din <= x"ff590485";
		wait for Clk_period;
		Addr <=  "00000011001101";
		Trees_din <= x"0afb1104";
		wait for Clk_period;
		Addr <=  "00000011001110";
		Trees_din <= x"00640485";
		wait for Clk_period;
		Addr <=  "00000011001111";
		Trees_din <= x"ff7b0485";
		wait for Clk_period;
		Addr <=  "00000011010000";
		Trees_din <= x"01fdd908";
		wait for Clk_period;
		Addr <=  "00000011010001";
		Trees_din <= x"11014304";
		wait for Clk_period;
		Addr <=  "00000011010010";
		Trees_din <= x"ffb70485";
		wait for Clk_period;
		Addr <=  "00000011010011";
		Trees_din <= x"013c0485";
		wait for Clk_period;
		Addr <=  "00000011010100";
		Trees_din <= x"0003aa04";
		wait for Clk_period;
		Addr <=  "00000011010101";
		Trees_din <= x"ff950485";
		wait for Clk_period;
		Addr <=  "00000011010110";
		Trees_din <= x"006e0485";
		wait for Clk_period;
		Addr <=  "00000011010111";
		Trees_din <= x"02094420";
		wait for Clk_period;
		Addr <=  "00000011011000";
		Trees_din <= x"010db610";
		wait for Clk_period;
		Addr <=  "00000011011001";
		Trees_din <= x"00090508";
		wait for Clk_period;
		Addr <=  "00000011011010";
		Trees_din <= x"0e009504";
		wait for Clk_period;
		Addr <=  "00000011011011";
		Trees_din <= x"00000485";
		wait for Clk_period;
		Addr <=  "00000011011100";
		Trees_din <= x"00a10485";
		wait for Clk_period;
		Addr <=  "00000011011101";
		Trees_din <= x"14006104";
		wait for Clk_period;
		Addr <=  "00000011011110";
		Trees_din <= x"00000485";
		wait for Clk_period;
		Addr <=  "00000011011111";
		Trees_din <= x"01070485";
		wait for Clk_period;
		Addr <=  "00000011100000";
		Trees_din <= x"12028708";
		wait for Clk_period;
		Addr <=  "00000011100001";
		Trees_din <= x"01107304";
		wait for Clk_period;
		Addr <=  "00000011100010";
		Trees_din <= x"ffd70485";
		wait for Clk_period;
		Addr <=  "00000011100011";
		Trees_din <= x"ff5c0485";
		wait for Clk_period;
		Addr <=  "00000011100100";
		Trees_din <= x"09004f04";
		wait for Clk_period;
		Addr <=  "00000011100101";
		Trees_din <= x"01a70485";
		wait for Clk_period;
		Addr <=  "00000011100110";
		Trees_din <= x"ffc90485";
		wait for Clk_period;
		Addr <=  "00000011100111";
		Trees_din <= x"17037310";
		wait for Clk_period;
		Addr <=  "00000011101000";
		Trees_din <= x"11007908";
		wait for Clk_period;
		Addr <=  "00000011101001";
		Trees_din <= x"1900a604";
		wait for Clk_period;
		Addr <=  "00000011101010";
		Trees_din <= x"ff7f0485";
		wait for Clk_period;
		Addr <=  "00000011101011";
		Trees_din <= x"00ac0485";
		wait for Clk_period;
		Addr <=  "00000011101100";
		Trees_din <= x"000b1e04";
		wait for Clk_period;
		Addr <=  "00000011101101";
		Trees_din <= x"ff5a0485";
		wait for Clk_period;
		Addr <=  "00000011101110";
		Trees_din <= x"ffc20485";
		wait for Clk_period;
		Addr <=  "00000011101111";
		Trees_din <= x"03facd04";
		wait for Clk_period;
		Addr <=  "00000011110000";
		Trees_din <= x"ff700485";
		wait for Clk_period;
		Addr <=  "00000011110001";
		Trees_din <= x"06f46304";
		wait for Clk_period;
		Addr <=  "00000011110010";
		Trees_din <= x"01840485";
		wait for Clk_period;
		Addr <=  "00000011110011";
		Trees_din <= x"00310485";
		wait for Clk_period;
		Addr <=  "00000011110100";
		Trees_din <= x"00100438";
		wait for Clk_period;
		Addr <=  "00000011110101";
		Trees_din <= x"010fff1c";
		wait for Clk_period;
		Addr <=  "00000011110110";
		Trees_din <= x"0208db0c";
		wait for Clk_period;
		Addr <=  "00000011110111";
		Trees_din <= x"12043608";
		wait for Clk_period;
		Addr <=  "00000011111000";
		Trees_din <= x"010a1f04";
		wait for Clk_period;
		Addr <=  "00000011111001";
		Trees_din <= x"01240485";
		wait for Clk_period;
		Addr <=  "00000011111010";
		Trees_din <= x"00a30485";
		wait for Clk_period;
		Addr <=  "00000011111011";
		Trees_din <= x"ff6c0485";
		wait for Clk_period;
		Addr <=  "00000011111100";
		Trees_din <= x"1402f408";
		wait for Clk_period;
		Addr <=  "00000011111101";
		Trees_din <= x"0d032a04";
		wait for Clk_period;
		Addr <=  "00000011111110";
		Trees_din <= x"ff920485";
		wait for Clk_period;
		Addr <=  "00000011111111";
		Trees_din <= x"008d0485";
		wait for Clk_period;
		Addr <=  "00000100000000";
		Trees_din <= x"03f82f04";
		wait for Clk_period;
		Addr <=  "00000100000001";
		Trees_din <= x"00420485";
		wait for Clk_period;
		Addr <=  "00000100000010";
		Trees_din <= x"01ae0485";
		wait for Clk_period;
		Addr <=  "00000100000011";
		Trees_din <= x"0a01d010";
		wait for Clk_period;
		Addr <=  "00000100000100";
		Trees_din <= x"05f9f308";
		wait for Clk_period;
		Addr <=  "00000100000101";
		Trees_din <= x"1a00f904";
		wait for Clk_period;
		Addr <=  "00000100000110";
		Trees_din <= x"ff5f0485";
		wait for Clk_period;
		Addr <=  "00000100000111";
		Trees_din <= x"003c0485";
		wait for Clk_period;
		Addr <=  "00000100001000";
		Trees_din <= x"07005704";
		wait for Clk_period;
		Addr <=  "00000100001001";
		Trees_din <= x"00d00485";
		wait for Clk_period;
		Addr <=  "00000100001010";
		Trees_din <= x"ffa20485";
		wait for Clk_period;
		Addr <=  "00000100001011";
		Trees_din <= x"03f84908";
		wait for Clk_period;
		Addr <=  "00000100001100";
		Trees_din <= x"0112d604";
		wait for Clk_period;
		Addr <=  "00000100001101";
		Trees_din <= x"01bd0485";
		wait for Clk_period;
		Addr <=  "00000100001110";
		Trees_din <= x"ffea0485";
		wait for Clk_period;
		Addr <=  "00000100001111";
		Trees_din <= x"ff750485";
		wait for Clk_period;
		Addr <=  "00000100010000";
		Trees_din <= x"0118031c";
		wait for Clk_period;
		Addr <=  "00000100010001";
		Trees_din <= x"00153210";
		wait for Clk_period;
		Addr <=  "00000100010010";
		Trees_din <= x"03f63f08";
		wait for Clk_period;
		Addr <=  "00000100010011";
		Trees_din <= x"09005b04";
		wait for Clk_period;
		Addr <=  "00000100010100";
		Trees_din <= x"00d70485";
		wait for Clk_period;
		Addr <=  "00000100010101";
		Trees_din <= x"ff8c0485";
		wait for Clk_period;
		Addr <=  "00000100010110";
		Trees_din <= x"1703f804";
		wait for Clk_period;
		Addr <=  "00000100010111";
		Trees_din <= x"01220485";
		wait for Clk_period;
		Addr <=  "00000100011000";
		Trees_din <= x"005c0485";
		wait for Clk_period;
		Addr <=  "00000100011001";
		Trees_din <= x"020d0604";
		wait for Clk_period;
		Addr <=  "00000100011010";
		Trees_din <= x"01300485";
		wait for Clk_period;
		Addr <=  "00000100011011";
		Trees_din <= x"00167604";
		wait for Clk_period;
		Addr <=  "00000100011100";
		Trees_din <= x"ff860485";
		wait for Clk_period;
		Addr <=  "00000100011101";
		Trees_din <= x"010d0485";
		wait for Clk_period;
		Addr <=  "00000100011110";
		Trees_din <= x"0d035304";
		wait for Clk_period;
		Addr <=  "00000100011111";
		Trees_din <= x"ff850485";
		wait for Clk_period;
		Addr <=  "00000100100000";
		Trees_din <= x"00340485";
		wait for Clk_period;
		Addr <=  "00000100100001";
		Trees_din <= x"0009b148";
		wait for Clk_period;
		Addr <=  "00000100100010";
		Trees_din <= x"0003aa20";
		wait for Clk_period;
		Addr <=  "00000100100011";
		Trees_din <= x"09003e08";
		wait for Clk_period;
		Addr <=  "00000100100100";
		Trees_din <= x"0f000704";
		wait for Clk_period;
		Addr <=  "00000100100101";
		Trees_din <= x"00ea0609";
		wait for Clk_period;
		Addr <=  "00000100100110";
		Trees_din <= x"ff8d0609";
		wait for Clk_period;
		Addr <=  "00000100100111";
		Trees_din <= x"1d005a10";
		wait for Clk_period;
		Addr <=  "00000100101000";
		Trees_din <= x"0000af08";
		wait for Clk_period;
		Addr <=  "00000100101001";
		Trees_din <= x"0803f904";
		wait for Clk_period;
		Addr <=  "00000100101010";
		Trees_din <= x"ff650609";
		wait for Clk_period;
		Addr <=  "00000100101011";
		Trees_din <= x"00300609";
		wait for Clk_period;
		Addr <=  "00000100101100";
		Trees_din <= x"0304d304";
		wait for Clk_period;
		Addr <=  "00000100101101";
		Trees_din <= x"ff770609";
		wait for Clk_period;
		Addr <=  "00000100101110";
		Trees_din <= x"00070609";
		wait for Clk_period;
		Addr <=  "00000100101111";
		Trees_din <= x"0d002a04";
		wait for Clk_period;
		Addr <=  "00000100110000";
		Trees_din <= x"01090609";
		wait for Clk_period;
		Addr <=  "00000100110001";
		Trees_din <= x"ff870609";
		wait for Clk_period;
		Addr <=  "00000100110010";
		Trees_din <= x"020b011c";
		wait for Clk_period;
		Addr <=  "00000100110011";
		Trees_din <= x"010f3710";
		wait for Clk_period;
		Addr <=  "00000100110100";
		Trees_din <= x"05fe9608";
		wait for Clk_period;
		Addr <=  "00000100110101";
		Trees_din <= x"01fec704";
		wait for Clk_period;
		Addr <=  "00000100110110";
		Trees_din <= x"00e90609";
		wait for Clk_period;
		Addr <=  "00000100110111";
		Trees_din <= x"00420609";
		wait for Clk_period;
		Addr <=  "00000100111000";
		Trees_din <= x"06fa5b04";
		wait for Clk_period;
		Addr <=  "00000100111001";
		Trees_din <= x"ff8d0609";
		wait for Clk_period;
		Addr <=  "00000100111010";
		Trees_din <= x"00a20609";
		wait for Clk_period;
		Addr <=  "00000100111011";
		Trees_din <= x"12028704";
		wait for Clk_period;
		Addr <=  "00000100111100";
		Trees_din <= x"ff630609";
		wait for Clk_period;
		Addr <=  "00000100111101";
		Trees_din <= x"14016404";
		wait for Clk_period;
		Addr <=  "00000100111110";
		Trees_din <= x"00f80609";
		wait for Clk_period;
		Addr <=  "00000100111111";
		Trees_din <= x"ff810609";
		wait for Clk_period;
		Addr <=  "00000101000000";
		Trees_din <= x"17036804";
		wait for Clk_period;
		Addr <=  "00000101000001";
		Trees_din <= x"ff600609";
		wait for Clk_period;
		Addr <=  "00000101000010";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00000101000011";
		Trees_din <= x"00d30609";
		wait for Clk_period;
		Addr <=  "00000101000100";
		Trees_din <= x"ff7b0609";
		wait for Clk_period;
		Addr <=  "00000101000101";
		Trees_din <= x"000f6f40";
		wait for Clk_period;
		Addr <=  "00000101000110";
		Trees_din <= x"0108f620";
		wait for Clk_period;
		Addr <=  "00000101000111";
		Trees_din <= x"02094410";
		wait for Clk_period;
		Addr <=  "00000101001000";
		Trees_din <= x"05024c08";
		wait for Clk_period;
		Addr <=  "00000101001001";
		Trees_din <= x"0b069b04";
		wait for Clk_period;
		Addr <=  "00000101001010";
		Trees_din <= x"00ec0609";
		wait for Clk_period;
		Addr <=  "00000101001011";
		Trees_din <= x"ffde0609";
		wait for Clk_period;
		Addr <=  "00000101001100";
		Trees_din <= x"13fe6804";
		wait for Clk_period;
		Addr <=  "00000101001101";
		Trees_din <= x"ff420609";
		wait for Clk_period;
		Addr <=  "00000101001110";
		Trees_din <= x"00400609";
		wait for Clk_period;
		Addr <=  "00000101001111";
		Trees_din <= x"0f022508";
		wait for Clk_period;
		Addr <=  "00000101010000";
		Trees_din <= x"1300b404";
		wait for Clk_period;
		Addr <=  "00000101010001";
		Trees_din <= x"ff7a0609";
		wait for Clk_period;
		Addr <=  "00000101010010";
		Trees_din <= x"00460609";
		wait for Clk_period;
		Addr <=  "00000101010011";
		Trees_din <= x"0afb1504";
		wait for Clk_period;
		Addr <=  "00000101010100";
		Trees_din <= x"01ac0609";
		wait for Clk_period;
		Addr <=  "00000101010101";
		Trees_din <= x"00100609";
		wait for Clk_period;
		Addr <=  "00000101010110";
		Trees_din <= x"0afc7c10";
		wait for Clk_period;
		Addr <=  "00000101010111";
		Trees_din <= x"05f9de08";
		wait for Clk_period;
		Addr <=  "00000101011000";
		Trees_din <= x"09005b04";
		wait for Clk_period;
		Addr <=  "00000101011001";
		Trees_din <= x"ff5b0609";
		wait for Clk_period;
		Addr <=  "00000101011010";
		Trees_din <= x"002d0609";
		wait for Clk_period;
		Addr <=  "00000101011011";
		Trees_din <= x"06f5ff04";
		wait for Clk_period;
		Addr <=  "00000101011100";
		Trees_din <= x"005e0609";
		wait for Clk_period;
		Addr <=  "00000101011101";
		Trees_din <= x"ff750609";
		wait for Clk_period;
		Addr <=  "00000101011110";
		Trees_din <= x"01139008";
		wait for Clk_period;
		Addr <=  "00000101011111";
		Trees_din <= x"10057a04";
		wait for Clk_period;
		Addr <=  "00000101100000";
		Trees_din <= x"00920609";
		wait for Clk_period;
		Addr <=  "00000101100001";
		Trees_din <= x"ff670609";
		wait for Clk_period;
		Addr <=  "00000101100010";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00000101100011";
		Trees_din <= x"00410609";
		wait for Clk_period;
		Addr <=  "00000101100100";
		Trees_din <= x"ff6e0609";
		wait for Clk_period;
		Addr <=  "00000101100101";
		Trees_din <= x"0111441c";
		wait for Clk_period;
		Addr <=  "00000101100110";
		Trees_din <= x"00153210";
		wait for Clk_period;
		Addr <=  "00000101100111";
		Trees_din <= x"01081408";
		wait for Clk_period;
		Addr <=  "00000101101000";
		Trees_din <= x"020e1a04";
		wait for Clk_period;
		Addr <=  "00000101101001";
		Trees_din <= x"00f10609";
		wait for Clk_period;
		Addr <=  "00000101101010";
		Trees_din <= x"00330609";
		wait for Clk_period;
		Addr <=  "00000101101011";
		Trees_din <= x"0c03c804";
		wait for Clk_period;
		Addr <=  "00000101101100";
		Trees_din <= x"00c90609";
		wait for Clk_period;
		Addr <=  "00000101101101";
		Trees_din <= x"00110609";
		wait for Clk_period;
		Addr <=  "00000101101110";
		Trees_din <= x"020d0604";
		wait for Clk_period;
		Addr <=  "00000101101111";
		Trees_din <= x"00f80609";
		wait for Clk_period;
		Addr <=  "00000101110000";
		Trees_din <= x"00167604";
		wait for Clk_period;
		Addr <=  "00000101110001";
		Trees_din <= x"ff8d0609";
		wait for Clk_period;
		Addr <=  "00000101110010";
		Trees_din <= x"00dd0609";
		wait for Clk_period;
		Addr <=  "00000101110011";
		Trees_din <= x"00167610";
		wait for Clk_period;
		Addr <=  "00000101110100";
		Trees_din <= x"0afcda08";
		wait for Clk_period;
		Addr <=  "00000101110101";
		Trees_din <= x"09005704";
		wait for Clk_period;
		Addr <=  "00000101110110";
		Trees_din <= x"ffb10609";
		wait for Clk_period;
		Addr <=  "00000101110111";
		Trees_din <= x"00830609";
		wait for Clk_period;
		Addr <=  "00000101111000";
		Trees_din <= x"0d016504";
		wait for Clk_period;
		Addr <=  "00000101111001";
		Trees_din <= x"00ea0609";
		wait for Clk_period;
		Addr <=  "00000101111010";
		Trees_din <= x"00160609";
		wait for Clk_period;
		Addr <=  "00000101111011";
		Trees_din <= x"1f000008";
		wait for Clk_period;
		Addr <=  "00000101111100";
		Trees_din <= x"10f74304";
		wait for Clk_period;
		Addr <=  "00000101111101";
		Trees_din <= x"00430609";
		wait for Clk_period;
		Addr <=  "00000101111110";
		Trees_din <= x"00fa0609";
		wait for Clk_period;
		Addr <=  "00000101111111";
		Trees_din <= x"01128f04";
		wait for Clk_period;
		Addr <=  "00000110000000";
		Trees_din <= x"00a20609";
		wait for Clk_period;
		Addr <=  "00000110000001";
		Trees_din <= x"ff650609";
		wait for Clk_period;
		Addr <=  "00000110000010";
		Trees_din <= x"000bca5c";
		wait for Clk_period;
		Addr <=  "00000110000011";
		Trees_din <= x"0003aa24";
		wait for Clk_period;
		Addr <=  "00000110000100";
		Trees_din <= x"09003e08";
		wait for Clk_period;
		Addr <=  "00000110000101";
		Trees_din <= x"0f000704";
		wait for Clk_period;
		Addr <=  "00000110000110";
		Trees_din <= x"00c10775";
		wait for Clk_period;
		Addr <=  "00000110000111";
		Trees_din <= x"ff950775";
		wait for Clk_period;
		Addr <=  "00000110001000";
		Trees_din <= x"0000af0c";
		wait for Clk_period;
		Addr <=  "00000110001001";
		Trees_din <= x"1204f608";
		wait for Clk_period;
		Addr <=  "00000110001010";
		Trees_din <= x"13f7ce04";
		wait for Clk_period;
		Addr <=  "00000110001011";
		Trees_din <= x"003b0775";
		wait for Clk_period;
		Addr <=  "00000110001100";
		Trees_din <= x"ff660775";
		wait for Clk_period;
		Addr <=  "00000110001101";
		Trees_din <= x"00430775";
		wait for Clk_period;
		Addr <=  "00000110001110";
		Trees_din <= x"01fdd908";
		wait for Clk_period;
		Addr <=  "00000110001111";
		Trees_din <= x"06f69704";
		wait for Clk_period;
		Addr <=  "00000110010000";
		Trees_din <= x"00c40775";
		wait for Clk_period;
		Addr <=  "00000110010001";
		Trees_din <= x"ffa80775";
		wait for Clk_period;
		Addr <=  "00000110010010";
		Trees_din <= x"0f000204";
		wait for Clk_period;
		Addr <=  "00000110010011";
		Trees_din <= x"00120775";
		wait for Clk_period;
		Addr <=  "00000110010100";
		Trees_din <= x"ff790775";
		wait for Clk_period;
		Addr <=  "00000110010101";
		Trees_din <= x"0209441c";
		wait for Clk_period;
		Addr <=  "00000110010110";
		Trees_din <= x"01092410";
		wait for Clk_period;
		Addr <=  "00000110010111";
		Trees_din <= x"06f55008";
		wait for Clk_period;
		Addr <=  "00000110011000";
		Trees_din <= x"11023204";
		wait for Clk_period;
		Addr <=  "00000110011001";
		Trees_din <= x"00660775";
		wait for Clk_period;
		Addr <=  "00000110011010";
		Trees_din <= x"01320775";
		wait for Clk_period;
		Addr <=  "00000110011011";
		Trees_din <= x"0f031504";
		wait for Clk_period;
		Addr <=  "00000110011100";
		Trees_din <= x"005d0775";
		wait for Clk_period;
		Addr <=  "00000110011101";
		Trees_din <= x"ffb10775";
		wait for Clk_period;
		Addr <=  "00000110011110";
		Trees_din <= x"0afb4d04";
		wait for Clk_period;
		Addr <=  "00000110011111";
		Trees_din <= x"ff5a0775";
		wait for Clk_period;
		Addr <=  "00000110100000";
		Trees_din <= x"09005d04";
		wait for Clk_period;
		Addr <=  "00000110100001";
		Trees_din <= x"00020775";
		wait for Clk_period;
		Addr <=  "00000110100010";
		Trees_din <= x"01590775";
		wait for Clk_period;
		Addr <=  "00000110100011";
		Trees_din <= x"17037310";
		wait for Clk_period;
		Addr <=  "00000110100100";
		Trees_din <= x"11007908";
		wait for Clk_period;
		Addr <=  "00000110100101";
		Trees_din <= x"1900a604";
		wait for Clk_period;
		Addr <=  "00000110100110";
		Trees_din <= x"ff8e0775";
		wait for Clk_period;
		Addr <=  "00000110100111";
		Trees_din <= x"00a40775";
		wait for Clk_period;
		Addr <=  "00000110101000";
		Trees_din <= x"01fdfc04";
		wait for Clk_period;
		Addr <=  "00000110101001";
		Trees_din <= x"ffd30775";
		wait for Clk_period;
		Addr <=  "00000110101010";
		Trees_din <= x"ff600775";
		wait for Clk_period;
		Addr <=  "00000110101011";
		Trees_din <= x"03facd04";
		wait for Clk_period;
		Addr <=  "00000110101100";
		Trees_din <= x"ff7b0775";
		wait for Clk_period;
		Addr <=  "00000110101101";
		Trees_din <= x"18004304";
		wait for Clk_period;
		Addr <=  "00000110101110";
		Trees_din <= x"01460775";
		wait for Clk_period;
		Addr <=  "00000110101111";
		Trees_din <= x"00290775";
		wait for Clk_period;
		Addr <=  "00000110110000";
		Trees_din <= x"00153238";
		wait for Clk_period;
		Addr <=  "00000110110001";
		Trees_din <= x"01139020";
		wait for Clk_period;
		Addr <=  "00000110110010";
		Trees_din <= x"02071410";
		wait for Clk_period;
		Addr <=  "00000110110011";
		Trees_din <= x"010a1f08";
		wait for Clk_period;
		Addr <=  "00000110110100";
		Trees_din <= x"16040004";
		wait for Clk_period;
		Addr <=  "00000110110101";
		Trees_din <= x"00c80775";
		wait for Clk_period;
		Addr <=  "00000110110110";
		Trees_din <= x"ffab0775";
		wait for Clk_period;
		Addr <=  "00000110110111";
		Trees_din <= x"0af78d04";
		wait for Clk_period;
		Addr <=  "00000110111000";
		Trees_din <= x"ff9f0775";
		wait for Clk_period;
		Addr <=  "00000110111001";
		Trees_din <= x"00930775";
		wait for Clk_period;
		Addr <=  "00000110111010";
		Trees_din <= x"11fdfc08";
		wait for Clk_period;
		Addr <=  "00000110111011";
		Trees_din <= x"0d00e504";
		wait for Clk_period;
		Addr <=  "00000110111100";
		Trees_din <= x"00970775";
		wait for Clk_period;
		Addr <=  "00000110111101";
		Trees_din <= x"ff5b0775";
		wait for Clk_period;
		Addr <=  "00000110111110";
		Trees_din <= x"0f000204";
		wait for Clk_period;
		Addr <=  "00000110111111";
		Trees_din <= x"ffe50775";
		wait for Clk_period;
		Addr <=  "00000111000000";
		Trees_din <= x"00880775";
		wait for Clk_period;
		Addr <=  "00000111000001";
		Trees_din <= x"12024c0c";
		wait for Clk_period;
		Addr <=  "00000111000010";
		Trees_din <= x"04fa9904";
		wait for Clk_period;
		Addr <=  "00000111000011";
		Trees_din <= x"ff600775";
		wait for Clk_period;
		Addr <=  "00000111000100";
		Trees_din <= x"00115704";
		wait for Clk_period;
		Addr <=  "00000111000101";
		Trees_din <= x"ff7d0775";
		wait for Clk_period;
		Addr <=  "00000111000110";
		Trees_din <= x"009b0775";
		wait for Clk_period;
		Addr <=  "00000111000111";
		Trees_din <= x"0bfb4404";
		wait for Clk_period;
		Addr <=  "00000111001000";
		Trees_din <= x"ff810775";
		wait for Clk_period;
		Addr <=  "00000111001001";
		Trees_din <= x"000f0704";
		wait for Clk_period;
		Addr <=  "00000111001010";
		Trees_din <= x"ffac0775";
		wait for Clk_period;
		Addr <=  "00000111001011";
		Trees_din <= x"00fd0775";
		wait for Clk_period;
		Addr <=  "00000111001100";
		Trees_din <= x"01128f0c";
		wait for Clk_period;
		Addr <=  "00000111001101";
		Trees_din <= x"020d0604";
		wait for Clk_period;
		Addr <=  "00000111001110";
		Trees_din <= x"00d80775";
		wait for Clk_period;
		Addr <=  "00000111001111";
		Trees_din <= x"00167604";
		wait for Clk_period;
		Addr <=  "00000111010000";
		Trees_din <= x"ff950775";
		wait for Clk_period;
		Addr <=  "00000111010001";
		Trees_din <= x"00bf0775";
		wait for Clk_period;
		Addr <=  "00000111010010";
		Trees_din <= x"01132a0c";
		wait for Clk_period;
		Addr <=  "00000111010011";
		Trees_din <= x"18004108";
		wait for Clk_period;
		Addr <=  "00000111010100";
		Trees_din <= x"00182604";
		wait for Clk_period;
		Addr <=  "00000111010101";
		Trees_din <= x"ffcd0775";
		wait for Clk_period;
		Addr <=  "00000111010110";
		Trees_din <= x"00c20775";
		wait for Clk_period;
		Addr <=  "00000111010111";
		Trees_din <= x"ff500775";
		wait for Clk_period;
		Addr <=  "00000111011000";
		Trees_din <= x"08032308";
		wait for Clk_period;
		Addr <=  "00000111011001";
		Trees_din <= x"1403eb04";
		wait for Clk_period;
		Addr <=  "00000111011010";
		Trees_din <= x"00d50775";
		wait for Clk_period;
		Addr <=  "00000111011011";
		Trees_din <= x"ffe40775";
		wait for Clk_period;
		Addr <=  "00000111011100";
		Trees_din <= x"ffde0775";
		wait for Clk_period;
		Addr <=  "00000111011101";
		Trees_din <= x"0009b148";
		wait for Clk_period;
		Addr <=  "00000111011110";
		Trees_din <= x"0003aa24";
		wait for Clk_period;
		Addr <=  "00000111011111";
		Trees_din <= x"1500760c";
		wait for Clk_period;
		Addr <=  "00000111100000";
		Trees_din <= x"0d002a08";
		wait for Clk_period;
		Addr <=  "00000111100001";
		Trees_din <= x"11026a04";
		wait for Clk_period;
		Addr <=  "00000111100010";
		Trees_din <= x"013408c9";
		wait for Clk_period;
		Addr <=  "00000111100011";
		Trees_din <= x"001808c9";
		wait for Clk_period;
		Addr <=  "00000111100100";
		Trees_din <= x"ff8308c9";
		wait for Clk_period;
		Addr <=  "00000111100101";
		Trees_din <= x"09003e08";
		wait for Clk_period;
		Addr <=  "00000111100110";
		Trees_din <= x"10043804";
		wait for Clk_period;
		Addr <=  "00000111100111";
		Trees_din <= x"00ae08c9";
		wait for Clk_period;
		Addr <=  "00000111101000";
		Trees_din <= x"ff9808c9";
		wait for Clk_period;
		Addr <=  "00000111101001";
		Trees_din <= x"0000af08";
		wait for Clk_period;
		Addr <=  "00000111101010";
		Trees_din <= x"1204f604";
		wait for Clk_period;
		Addr <=  "00000111101011";
		Trees_din <= x"ff6b08c9";
		wait for Clk_period;
		Addr <=  "00000111101100";
		Trees_din <= x"004108c9";
		wait for Clk_period;
		Addr <=  "00000111101101";
		Trees_din <= x"0bf94004";
		wait for Clk_period;
		Addr <=  "00000111101110";
		Trees_din <= x"006d08c9";
		wait for Clk_period;
		Addr <=  "00000111101111";
		Trees_din <= x"ff9608c9";
		wait for Clk_period;
		Addr <=  "00000111110000";
		Trees_din <= x"020cbe20";
		wait for Clk_period;
		Addr <=  "00000111110001";
		Trees_din <= x"16015b10";
		wait for Clk_period;
		Addr <=  "00000111110010";
		Trees_din <= x"1201e208";
		wait for Clk_period;
		Addr <=  "00000111110011";
		Trees_din <= x"0af7dc04";
		wait for Clk_period;
		Addr <=  "00000111110100";
		Trees_din <= x"008408c9";
		wait for Clk_period;
		Addr <=  "00000111110101";
		Trees_din <= x"ff5808c9";
		wait for Clk_period;
		Addr <=  "00000111110110";
		Trees_din <= x"1b003804";
		wait for Clk_period;
		Addr <=  "00000111110111";
		Trees_din <= x"ffa608c9";
		wait for Clk_period;
		Addr <=  "00000111111000";
		Trees_din <= x"007508c9";
		wait for Clk_period;
		Addr <=  "00000111111001";
		Trees_din <= x"18003d08";
		wait for Clk_period;
		Addr <=  "00000111111010";
		Trees_din <= x"07005604";
		wait for Clk_period;
		Addr <=  "00000111111011";
		Trees_din <= x"002208c9";
		wait for Clk_period;
		Addr <=  "00000111111100";
		Trees_din <= x"ff5608c9";
		wait for Clk_period;
		Addr <=  "00000111111101";
		Trees_din <= x"04fc5b04";
		wait for Clk_period;
		Addr <=  "00000111111110";
		Trees_din <= x"ffdc08c9";
		wait for Clk_period;
		Addr <=  "00000111111111";
		Trees_din <= x"008f08c9";
		wait for Clk_period;
		Addr <=  "00001000000000";
		Trees_din <= x"ff6708c9";
		wait for Clk_period;
		Addr <=  "00001000000001";
		Trees_din <= x"0015323c";
		wait for Clk_period;
		Addr <=  "00001000000010";
		Trees_din <= x"0108bd20";
		wait for Clk_period;
		Addr <=  "00001000000011";
		Trees_din <= x"020abe10";
		wait for Clk_period;
		Addr <=  "00001000000100";
		Trees_din <= x"05034408";
		wait for Clk_period;
		Addr <=  "00001000000101";
		Trees_din <= x"07006004";
		wait for Clk_period;
		Addr <=  "00001000000110";
		Trees_din <= x"00ab08c9";
		wait for Clk_period;
		Addr <=  "00001000000111";
		Trees_din <= x"ffa008c9";
		wait for Clk_period;
		Addr <=  "00001000001000";
		Trees_din <= x"16003904";
		wait for Clk_period;
		Addr <=  "00001000001001";
		Trees_din <= x"ff4808c9";
		wait for Clk_period;
		Addr <=  "00001000001010";
		Trees_din <= x"004908c9";
		wait for Clk_period;
		Addr <=  "00001000001011";
		Trees_din <= x"000f0708";
		wait for Clk_period;
		Addr <=  "00001000001100";
		Trees_din <= x"11007904";
		wait for Clk_period;
		Addr <=  "00001000001101";
		Trees_din <= x"00b708c9";
		wait for Clk_period;
		Addr <=  "00001000001110";
		Trees_din <= x"ff9c08c9";
		wait for Clk_period;
		Addr <=  "00001000001111";
		Trees_din <= x"17007d04";
		wait for Clk_period;
		Addr <=  "00001000010000";
		Trees_din <= x"00c808c9";
		wait for Clk_period;
		Addr <=  "00001000010001";
		Trees_din <= x"000208c9";
		wait for Clk_period;
		Addr <=  "00001000010010";
		Trees_din <= x"0113e910";
		wait for Clk_period;
		Addr <=  "00001000010011";
		Trees_din <= x"000d2308";
		wait for Clk_period;
		Addr <=  "00001000010100";
		Trees_din <= x"0f03f604";
		wait for Clk_period;
		Addr <=  "00001000010101";
		Trees_din <= x"fffd08c9";
		wait for Clk_period;
		Addr <=  "00001000010110";
		Trees_din <= x"013208c9";
		wait for Clk_period;
		Addr <=  "00001000010111";
		Trees_din <= x"06f35804";
		wait for Clk_period;
		Addr <=  "00001000011000";
		Trees_din <= x"00c008c9";
		wait for Clk_period;
		Addr <=  "00001000011001";
		Trees_din <= x"006108c9";
		wait for Clk_period;
		Addr <=  "00001000011010";
		Trees_din <= x"0efa8a04";
		wait for Clk_period;
		Addr <=  "00001000011011";
		Trees_din <= x"00a908c9";
		wait for Clk_period;
		Addr <=  "00001000011100";
		Trees_din <= x"0011ff04";
		wait for Clk_period;
		Addr <=  "00001000011101";
		Trees_din <= x"ff6608c9";
		wait for Clk_period;
		Addr <=  "00001000011110";
		Trees_din <= x"001b08c9";
		wait for Clk_period;
		Addr <=  "00001000011111";
		Trees_din <= x"010d4f14";
		wait for Clk_period;
		Addr <=  "00001000100000";
		Trees_din <= x"020d060c";
		wait for Clk_period;
		Addr <=  "00001000100001";
		Trees_din <= x"1a013704";
		wait for Clk_period;
		Addr <=  "00001000100010";
		Trees_din <= x"00c508c9";
		wait for Clk_period;
		Addr <=  "00001000100011";
		Trees_din <= x"0bfb4404";
		wait for Clk_period;
		Addr <=  "00001000100100";
		Trees_din <= x"ffe508c9";
		wait for Clk_period;
		Addr <=  "00001000100101";
		Trees_din <= x"009908c9";
		wait for Clk_period;
		Addr <=  "00001000100110";
		Trees_din <= x"00167604";
		wait for Clk_period;
		Addr <=  "00001000100111";
		Trees_din <= x"ff9c08c9";
		wait for Clk_period;
		Addr <=  "00001000101000";
		Trees_din <= x"009f08c9";
		wait for Clk_period;
		Addr <=  "00001000101001";
		Trees_din <= x"0bf88604";
		wait for Clk_period;
		Addr <=  "00001000101010";
		Trees_din <= x"ffa708c9";
		wait for Clk_period;
		Addr <=  "00001000101011";
		Trees_din <= x"03f7b308";
		wait for Clk_period;
		Addr <=  "00001000101100";
		Trees_din <= x"00167604";
		wait for Clk_period;
		Addr <=  "00001000101101";
		Trees_din <= x"006408c9";
		wait for Clk_period;
		Addr <=  "00001000101110";
		Trees_din <= x"00b508c9";
		wait for Clk_period;
		Addr <=  "00001000101111";
		Trees_din <= x"08022004";
		wait for Clk_period;
		Addr <=  "00001000110000";
		Trees_din <= x"ff6008c9";
		wait for Clk_period;
		Addr <=  "00001000110001";
		Trees_din <= x"007008c9";
		wait for Clk_period;
		Addr <=  "00001000110010";
		Trees_din <= x"000ceb70";
		wait for Clk_period;
		Addr <=  "00001000110011";
		Trees_din <= x"00058434";
		wait for Clk_period;
		Addr <=  "00001000110100";
		Trees_din <= x"0000af18";
		wait for Clk_period;
		Addr <=  "00001000110101";
		Trees_din <= x"1a010510";
		wait for Clk_period;
		Addr <=  "00001000110110";
		Trees_din <= x"1703f208";
		wait for Clk_period;
		Addr <=  "00001000110111";
		Trees_din <= x"1204f604";
		wait for Clk_period;
		Addr <=  "00001000111000";
		Trees_din <= x"ff660a55";
		wait for Clk_period;
		Addr <=  "00001000111001";
		Trees_din <= x"00400a55";
		wait for Clk_period;
		Addr <=  "00001000111010";
		Trees_din <= x"04fe3404";
		wait for Clk_period;
		Addr <=  "00001000111011";
		Trees_din <= x"00c10a55";
		wait for Clk_period;
		Addr <=  "00001000111100";
		Trees_din <= x"ff8b0a55";
		wait for Clk_period;
		Addr <=  "00001000111101";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00001000111110";
		Trees_din <= x"00ca0a55";
		wait for Clk_period;
		Addr <=  "00001000111111";
		Trees_din <= x"ff8c0a55";
		wait for Clk_period;
		Addr <=  "00001001000000";
		Trees_din <= x"03fd840c";
		wait for Clk_period;
		Addr <=  "00001001000001";
		Trees_din <= x"06091b08";
		wait for Clk_period;
		Addr <=  "00001001000010";
		Trees_din <= x"22000004";
		wait for Clk_period;
		Addr <=  "00001001000011";
		Trees_din <= x"ff610a55";
		wait for Clk_period;
		Addr <=  "00001001000100";
		Trees_din <= x"00350a55";
		wait for Clk_period;
		Addr <=  "00001001000101";
		Trees_din <= x"003b0a55";
		wait for Clk_period;
		Addr <=  "00001001000110";
		Trees_din <= x"1603fe08";
		wait for Clk_period;
		Addr <=  "00001001000111";
		Trees_din <= x"07005804";
		wait for Clk_period;
		Addr <=  "00001001001000";
		Trees_din <= x"001c0a55";
		wait for Clk_period;
		Addr <=  "00001001001001";
		Trees_din <= x"ff950a55";
		wait for Clk_period;
		Addr <=  "00001001001010";
		Trees_din <= x"1003b904";
		wait for Clk_period;
		Addr <=  "00001001001011";
		Trees_din <= x"01690a55";
		wait for Clk_period;
		Addr <=  "00001001001100";
		Trees_din <= x"00460a55";
		wait for Clk_period;
		Addr <=  "00001001001101";
		Trees_din <= x"03fa8720";
		wait for Clk_period;
		Addr <=  "00001001001110";
		Trees_din <= x"08025910";
		wait for Clk_period;
		Addr <=  "00001001001111";
		Trees_din <= x"1a00d108";
		wait for Clk_period;
		Addr <=  "00001001010000";
		Trees_din <= x"1a00b204";
		wait for Clk_period;
		Addr <=  "00001001010001";
		Trees_din <= x"ff900a55";
		wait for Clk_period;
		Addr <=  "00001001010010";
		Trees_din <= x"002f0a55";
		wait for Clk_period;
		Addr <=  "00001001010011";
		Trees_din <= x"0d038804";
		wait for Clk_period;
		Addr <=  "00001001010100";
		Trees_din <= x"ff5e0a55";
		wait for Clk_period;
		Addr <=  "00001001010101";
		Trees_din <= x"00230a55";
		wait for Clk_period;
		Addr <=  "00001001010110";
		Trees_din <= x"0c01f408";
		wait for Clk_period;
		Addr <=  "00001001010111";
		Trees_din <= x"18004404";
		wait for Clk_period;
		Addr <=  "00001001011000";
		Trees_din <= x"01340a55";
		wait for Clk_period;
		Addr <=  "00001001011001";
		Trees_din <= x"ff9d0a55";
		wait for Clk_period;
		Addr <=  "00001001011010";
		Trees_din <= x"05fba104";
		wait for Clk_period;
		Addr <=  "00001001011011";
		Trees_din <= x"ff720a55";
		wait for Clk_period;
		Addr <=  "00001001011100";
		Trees_din <= x"00230a55";
		wait for Clk_period;
		Addr <=  "00001001011101";
		Trees_din <= x"09005810";
		wait for Clk_period;
		Addr <=  "00001001011110";
		Trees_din <= x"01020f08";
		wait for Clk_period;
		Addr <=  "00001001011111";
		Trees_din <= x"0afcc204";
		wait for Clk_period;
		Addr <=  "00001001100000";
		Trees_din <= x"00d70a55";
		wait for Clk_period;
		Addr <=  "00001001100001";
		Trees_din <= x"00240a55";
		wait for Clk_period;
		Addr <=  "00001001100010";
		Trees_din <= x"04fd7904";
		wait for Clk_period;
		Addr <=  "00001001100011";
		Trees_din <= x"ff850a55";
		wait for Clk_period;
		Addr <=  "00001001100100";
		Trees_din <= x"00450a55";
		wait for Clk_period;
		Addr <=  "00001001100101";
		Trees_din <= x"0b055908";
		wait for Clk_period;
		Addr <=  "00001001100110";
		Trees_din <= x"0afb1e04";
		wait for Clk_period;
		Addr <=  "00001001100111";
		Trees_din <= x"fff00a55";
		wait for Clk_period;
		Addr <=  "00001001101000";
		Trees_din <= x"00d60a55";
		wait for Clk_period;
		Addr <=  "00001001101001";
		Trees_din <= x"ff710a55";
		wait for Clk_period;
		Addr <=  "00001001101010";
		Trees_din <= x"0016763c";
		wait for Clk_period;
		Addr <=  "00001001101011";
		Trees_din <= x"01082a20";
		wait for Clk_period;
		Addr <=  "00001001101100";
		Trees_din <= x"0205a110";
		wait for Clk_period;
		Addr <=  "00001001101101";
		Trees_din <= x"11fb6308";
		wait for Clk_period;
		Addr <=  "00001001101110";
		Trees_din <= x"0f014e04";
		wait for Clk_period;
		Addr <=  "00001001101111";
		Trees_din <= x"ff720a55";
		wait for Clk_period;
		Addr <=  "00001001110000";
		Trees_din <= x"007b0a55";
		wait for Clk_period;
		Addr <=  "00001001110001";
		Trees_din <= x"0501a404";
		wait for Clk_period;
		Addr <=  "00001001110010";
		Trees_din <= x"00ac0a55";
		wait for Clk_period;
		Addr <=  "00001001110011";
		Trees_din <= x"00510a55";
		wait for Clk_period;
		Addr <=  "00001001110100";
		Trees_din <= x"0b028808";
		wait for Clk_period;
		Addr <=  "00001001110101";
		Trees_din <= x"020e8d04";
		wait for Clk_period;
		Addr <=  "00001001110110";
		Trees_din <= x"00a50a55";
		wait for Clk_period;
		Addr <=  "00001001110111";
		Trees_din <= x"ffc40a55";
		wait for Clk_period;
		Addr <=  "00001001111000";
		Trees_din <= x"17000004";
		wait for Clk_period;
		Addr <=  "00001001111001";
		Trees_din <= x"ff790a55";
		wait for Clk_period;
		Addr <=  "00001001111010";
		Trees_din <= x"00530a55";
		wait for Clk_period;
		Addr <=  "00001001111011";
		Trees_din <= x"0c03c80c";
		wait for Clk_period;
		Addr <=  "00001001111100";
		Trees_din <= x"01173e08";
		wait for Clk_period;
		Addr <=  "00001001111101";
		Trees_din <= x"07005b04";
		wait for Clk_period;
		Addr <=  "00001001111110";
		Trees_din <= x"006f0a55";
		wait for Clk_period;
		Addr <=  "00001001111111";
		Trees_din <= x"00120a55";
		wait for Clk_period;
		Addr <=  "00001010000000";
		Trees_din <= x"ff7c0a55";
		wait for Clk_period;
		Addr <=  "00001010000001";
		Trees_din <= x"0c03dd08";
		wait for Clk_period;
		Addr <=  "00001010000010";
		Trees_din <= x"0f002c04";
		wait for Clk_period;
		Addr <=  "00001010000011";
		Trees_din <= x"00070a55";
		wait for Clk_period;
		Addr <=  "00001010000100";
		Trees_din <= x"ff190a55";
		wait for Clk_period;
		Addr <=  "00001010000101";
		Trees_din <= x"03f74704";
		wait for Clk_period;
		Addr <=  "00001010000110";
		Trees_din <= x"00c60a55";
		wait for Clk_period;
		Addr <=  "00001010000111";
		Trees_din <= x"ffc90a55";
		wait for Clk_period;
		Addr <=  "00001010001000";
		Trees_din <= x"01164210";
		wait for Clk_period;
		Addr <=  "00001010001001";
		Trees_din <= x"010d4f04";
		wait for Clk_period;
		Addr <=  "00001010001010";
		Trees_din <= x"00b80a55";
		wait for Clk_period;
		Addr <=  "00001010001011";
		Trees_din <= x"0bf88604";
		wait for Clk_period;
		Addr <=  "00001010001100";
		Trees_din <= x"ffa40a55";
		wait for Clk_period;
		Addr <=  "00001010001101";
		Trees_din <= x"03f7b304";
		wait for Clk_period;
		Addr <=  "00001010001110";
		Trees_din <= x"00a70a55";
		wait for Clk_period;
		Addr <=  "00001010001111";
		Trees_din <= x"ffd90a55";
		wait for Clk_period;
		Addr <=  "00001010010000";
		Trees_din <= x"0b039108";
		wait for Clk_period;
		Addr <=  "00001010010001";
		Trees_din <= x"09005204";
		wait for Clk_period;
		Addr <=  "00001010010010";
		Trees_din <= x"00140a55";
		wait for Clk_period;
		Addr <=  "00001010010011";
		Trees_din <= x"ff8e0a55";
		wait for Clk_period;
		Addr <=  "00001010010100";
		Trees_din <= x"00950a55";
		wait for Clk_period;
		Addr <=  "00001010010101";
		Trees_din <= x"000f6f64";
		wait for Clk_period;
		Addr <=  "00001010010110";
		Trees_din <= x"0004a13c";
		wait for Clk_period;
		Addr <=  "00001010010111";
		Trees_din <= x"0000af1c";
		wait for Clk_period;
		Addr <=  "00001010011000";
		Trees_din <= x"1a010510";
		wait for Clk_period;
		Addr <=  "00001010011001";
		Trees_din <= x"1703f208";
		wait for Clk_period;
		Addr <=  "00001010011010";
		Trees_din <= x"1204f604";
		wait for Clk_period;
		Addr <=  "00001010011011";
		Trees_din <= x"ff690bd9";
		wait for Clk_period;
		Addr <=  "00001010011100";
		Trees_din <= x"003e0bd9";
		wait for Clk_period;
		Addr <=  "00001010011101";
		Trees_din <= x"06f8e004";
		wait for Clk_period;
		Addr <=  "00001010011110";
		Trees_din <= x"ff910bd9";
		wait for Clk_period;
		Addr <=  "00001010011111";
		Trees_din <= x"00b60bd9";
		wait for Clk_period;
		Addr <=  "00001010100000";
		Trees_din <= x"20040008";
		wait for Clk_period;
		Addr <=  "00001010100001";
		Trees_din <= x"06f81604";
		wait for Clk_period;
		Addr <=  "00001010100010";
		Trees_din <= x"00d30bd9";
		wait for Clk_period;
		Addr <=  "00001010100011";
		Trees_din <= x"00300bd9";
		wait for Clk_period;
		Addr <=  "00001010100100";
		Trees_din <= x"ff930bd9";
		wait for Clk_period;
		Addr <=  "00001010100101";
		Trees_din <= x"04025d10";
		wait for Clk_period;
		Addr <=  "00001010100110";
		Trees_din <= x"0d03ae08";
		wait for Clk_period;
		Addr <=  "00001010100111";
		Trees_din <= x"0ef9a204";
		wait for Clk_period;
		Addr <=  "00001010101000";
		Trees_din <= x"000b0bd9";
		wait for Clk_period;
		Addr <=  "00001010101001";
		Trees_din <= x"ff610bd9";
		wait for Clk_period;
		Addr <=  "00001010101010";
		Trees_din <= x"07005704";
		wait for Clk_period;
		Addr <=  "00001010101011";
		Trees_din <= x"00ab0bd9";
		wait for Clk_period;
		Addr <=  "00001010101100";
		Trees_din <= x"ff8e0bd9";
		wait for Clk_period;
		Addr <=  "00001010101101";
		Trees_din <= x"08021408";
		wait for Clk_period;
		Addr <=  "00001010101110";
		Trees_din <= x"18004a04";
		wait for Clk_period;
		Addr <=  "00001010101111";
		Trees_din <= x"ffac0bd9";
		wait for Clk_period;
		Addr <=  "00001010110000";
		Trees_din <= x"00710bd9";
		wait for Clk_period;
		Addr <=  "00001010110001";
		Trees_din <= x"08029604";
		wait for Clk_period;
		Addr <=  "00001010110010";
		Trees_din <= x"01460bd9";
		wait for Clk_period;
		Addr <=  "00001010110011";
		Trees_din <= x"ffc20bd9";
		wait for Clk_period;
		Addr <=  "00001010110100";
		Trees_din <= x"03f5ed08";
		wait for Clk_period;
		Addr <=  "00001010110101";
		Trees_din <= x"000f0704";
		wait for Clk_period;
		Addr <=  "00001010110110";
		Trees_din <= x"ff620bd9";
		wait for Clk_period;
		Addr <=  "00001010110111";
		Trees_din <= x"00490bd9";
		wait for Clk_period;
		Addr <=  "00001010111000";
		Trees_din <= x"0101df10";
		wait for Clk_period;
		Addr <=  "00001010111001";
		Trees_din <= x"05011d08";
		wait for Clk_period;
		Addr <=  "00001010111010";
		Trees_din <= x"0afcad04";
		wait for Clk_period;
		Addr <=  "00001010111011";
		Trees_din <= x"00ba0bd9";
		wait for Clk_period;
		Addr <=  "00001010111100";
		Trees_din <= x"004a0bd9";
		wait for Clk_period;
		Addr <=  "00001010111101";
		Trees_din <= x"11045104";
		wait for Clk_period;
		Addr <=  "00001010111110";
		Trees_din <= x"ff6b0bd9";
		wait for Clk_period;
		Addr <=  "00001010111111";
		Trees_din <= x"009a0bd9";
		wait for Clk_period;
		Addr <=  "00001011000000";
		Trees_din <= x"06f75208";
		wait for Clk_period;
		Addr <=  "00001011000001";
		Trees_din <= x"10059704";
		wait for Clk_period;
		Addr <=  "00001011000010";
		Trees_din <= x"00470bd9";
		wait for Clk_period;
		Addr <=  "00001011000011";
		Trees_din <= x"ff8c0bd9";
		wait for Clk_period;
		Addr <=  "00001011000100";
		Trees_din <= x"09005804";
		wait for Clk_period;
		Addr <=  "00001011000101";
		Trees_din <= x"ffbd0bd9";
		wait for Clk_period;
		Addr <=  "00001011000110";
		Trees_din <= x"00730bd9";
		wait for Clk_period;
		Addr <=  "00001011000111";
		Trees_din <= x"00167640";
		wait for Clk_period;
		Addr <=  "00001011001000";
		Trees_din <= x"010d4f20";
		wait for Clk_period;
		Addr <=  "00001011001001";
		Trees_din <= x"0c019510";
		wait for Clk_period;
		Addr <=  "00001011001010";
		Trees_din <= x"0d003408";
		wait for Clk_period;
		Addr <=  "00001011001011";
		Trees_din <= x"01096904";
		wait for Clk_period;
		Addr <=  "00001011001100";
		Trees_din <= x"00970bd9";
		wait for Clk_period;
		Addr <=  "00001011001101";
		Trees_din <= x"fffe0bd9";
		wait for Clk_period;
		Addr <=  "00001011001110";
		Trees_din <= x"0b059404";
		wait for Clk_period;
		Addr <=  "00001011001111";
		Trees_din <= x"00b60bd9";
		wait for Clk_period;
		Addr <=  "00001011010000";
		Trees_din <= x"000a0bd9";
		wait for Clk_period;
		Addr <=  "00001011010001";
		Trees_din <= x"02097608";
		wait for Clk_period;
		Addr <=  "00001011010010";
		Trees_din <= x"1b003a04";
		wait for Clk_period;
		Addr <=  "00001011010011";
		Trees_din <= x"00570bd9";
		wait for Clk_period;
		Addr <=  "00001011010100";
		Trees_din <= x"00980bd9";
		wait for Clk_period;
		Addr <=  "00001011010101";
		Trees_din <= x"06f4d304";
		wait for Clk_period;
		Addr <=  "00001011010110";
		Trees_din <= x"00700bd9";
		wait for Clk_period;
		Addr <=  "00001011010111";
		Trees_din <= x"ff6a0bd9";
		wait for Clk_period;
		Addr <=  "00001011011000";
		Trees_din <= x"1d004110";
		wait for Clk_period;
		Addr <=  "00001011011001";
		Trees_din <= x"0c02d908";
		wait for Clk_period;
		Addr <=  "00001011011010";
		Trees_din <= x"0015c504";
		wait for Clk_period;
		Addr <=  "00001011011011";
		Trees_din <= x"00b00bd9";
		wait for Clk_period;
		Addr <=  "00001011011100";
		Trees_din <= x"ffe20bd9";
		wait for Clk_period;
		Addr <=  "00001011011101";
		Trees_din <= x"0802f004";
		wait for Clk_period;
		Addr <=  "00001011011110";
		Trees_din <= x"003d0bd9";
		wait for Clk_period;
		Addr <=  "00001011011111";
		Trees_din <= x"ff3c0bd9";
		wait for Clk_period;
		Addr <=  "00001011100000";
		Trees_din <= x"19008608";
		wait for Clk_period;
		Addr <=  "00001011100001";
		Trees_din <= x"01139004";
		wait for Clk_period;
		Addr <=  "00001011100010";
		Trees_din <= x"00a50bd9";
		wait for Clk_period;
		Addr <=  "00001011100011";
		Trees_din <= x"fff20bd9";
		wait for Clk_period;
		Addr <=  "00001011100100";
		Trees_din <= x"21000004";
		wait for Clk_period;
		Addr <=  "00001011100101";
		Trees_din <= x"ffd00bd9";
		wait for Clk_period;
		Addr <=  "00001011100110";
		Trees_din <= x"00bf0bd9";
		wait for Clk_period;
		Addr <=  "00001011100111";
		Trees_din <= x"010d4f0c";
		wait for Clk_period;
		Addr <=  "00001011101000";
		Trees_din <= x"0a07cb04";
		wait for Clk_period;
		Addr <=  "00001011101001";
		Trees_din <= x"00af0bd9";
		wait for Clk_period;
		Addr <=  "00001011101010";
		Trees_din <= x"15009404";
		wait for Clk_period;
		Addr <=  "00001011101011";
		Trees_din <= x"ffc40bd9";
		wait for Clk_period;
		Addr <=  "00001011101100";
		Trees_din <= x"008a0bd9";
		wait for Clk_period;
		Addr <=  "00001011101101";
		Trees_din <= x"0bf88604";
		wait for Clk_period;
		Addr <=  "00001011101110";
		Trees_din <= x"ffa70bd9";
		wait for Clk_period;
		Addr <=  "00001011101111";
		Trees_din <= x"03f7b308";
		wait for Clk_period;
		Addr <=  "00001011110000";
		Trees_din <= x"0a079004";
		wait for Clk_period;
		Addr <=  "00001011110001";
		Trees_din <= x"00970bd9";
		wait for Clk_period;
		Addr <=  "00001011110010";
		Trees_din <= x"fff00bd9";
		wait for Clk_period;
		Addr <=  "00001011110011";
		Trees_din <= x"00170d04";
		wait for Clk_period;
		Addr <=  "00001011110100";
		Trees_din <= x"00640bd9";
		wait for Clk_period;
		Addr <=  "00001011110101";
		Trees_din <= x"ff600bd9";
		wait for Clk_period;
		Addr <=  "00001011110110";
		Trees_din <= x"00119270";
		wait for Clk_period;
		Addr <=  "00001011110111";
		Trees_din <= x"00079034";
		wait for Clk_period;
		Addr <=  "00001011111000";
		Trees_din <= x"0000af18";
		wait for Clk_period;
		Addr <=  "00001011111001";
		Trees_din <= x"02fba50c";
		wait for Clk_period;
		Addr <=  "00001011111010";
		Trees_din <= x"14003304";
		wait for Clk_period;
		Addr <=  "00001011111011";
		Trees_din <= x"00f40d65";
		wait for Clk_period;
		Addr <=  "00001011111100";
		Trees_din <= x"1e005604";
		wait for Clk_period;
		Addr <=  "00001011111101";
		Trees_din <= x"002c0d65";
		wait for Clk_period;
		Addr <=  "00001011111110";
		Trees_din <= x"ff850d65";
		wait for Clk_period;
		Addr <=  "00001011111111";
		Trees_din <= x"1204f608";
		wait for Clk_period;
		Addr <=  "00001100000000";
		Trees_din <= x"18003104";
		wait for Clk_period;
		Addr <=  "00001100000001";
		Trees_din <= x"001c0d65";
		wait for Clk_period;
		Addr <=  "00001100000010";
		Trees_din <= x"ff6b0d65";
		wait for Clk_period;
		Addr <=  "00001100000011";
		Trees_din <= x"00390d65";
		wait for Clk_period;
		Addr <=  "00001100000100";
		Trees_din <= x"01fdeb0c";
		wait for Clk_period;
		Addr <=  "00001100000101";
		Trees_din <= x"11fed304";
		wait for Clk_period;
		Addr <=  "00001100000110";
		Trees_din <= x"ff760d65";
		wait for Clk_period;
		Addr <=  "00001100000111";
		Trees_din <= x"06f69704";
		wait for Clk_period;
		Addr <=  "00001100001000";
		Trees_din <= x"00bb0d65";
		wait for Clk_period;
		Addr <=  "00001100001001";
		Trees_din <= x"001c0d65";
		wait for Clk_period;
		Addr <=  "00001100001010";
		Trees_din <= x"0e01f008";
		wait for Clk_period;
		Addr <=  "00001100001011";
		Trees_din <= x"09005404";
		wait for Clk_period;
		Addr <=  "00001100001100";
		Trees_din <= x"ff7d0d65";
		wait for Clk_period;
		Addr <=  "00001100001101";
		Trees_din <= x"ffde0d65";
		wait for Clk_period;
		Addr <=  "00001100001110";
		Trees_din <= x"03fce704";
		wait for Clk_period;
		Addr <=  "00001100001111";
		Trees_din <= x"ff7e0d65";
		wait for Clk_period;
		Addr <=  "00001100010000";
		Trees_din <= x"00440d65";
		wait for Clk_period;
		Addr <=  "00001100010001";
		Trees_din <= x"04fc431c";
		wait for Clk_period;
		Addr <=  "00001100010010";
		Trees_din <= x"0009b10c";
		wait for Clk_period;
		Addr <=  "00001100010011";
		Trees_din <= x"10f7fb04";
		wait for Clk_period;
		Addr <=  "00001100010100";
		Trees_din <= x"008a0d65";
		wait for Clk_period;
		Addr <=  "00001100010101";
		Trees_din <= x"1d003804";
		wait for Clk_period;
		Addr <=  "00001100010110";
		Trees_din <= x"003c0d65";
		wait for Clk_period;
		Addr <=  "00001100010111";
		Trees_din <= x"ff710d65";
		wait for Clk_period;
		Addr <=  "00001100011000";
		Trees_din <= x"1f000008";
		wait for Clk_period;
		Addr <=  "00001100011001";
		Trees_din <= x"08001504";
		wait for Clk_period;
		Addr <=  "00001100011010";
		Trees_din <= x"006f0d65";
		wait for Clk_period;
		Addr <=  "00001100011011";
		Trees_din <= x"00000d65";
		wait for Clk_period;
		Addr <=  "00001100011100";
		Trees_din <= x"03f55804";
		wait for Clk_period;
		Addr <=  "00001100011101";
		Trees_din <= x"ff7f0d65";
		wait for Clk_period;
		Addr <=  "00001100011110";
		Trees_din <= x"00ab0d65";
		wait for Clk_period;
		Addr <=  "00001100011111";
		Trees_din <= x"09005810";
		wait for Clk_period;
		Addr <=  "00001100100000";
		Trees_din <= x"000d2308";
		wait for Clk_period;
		Addr <=  "00001100100001";
		Trees_din <= x"04fea404";
		wait for Clk_period;
		Addr <=  "00001100100010";
		Trees_din <= x"ffd80d65";
		wait for Clk_period;
		Addr <=  "00001100100011";
		Trees_din <= x"00460d65";
		wait for Clk_period;
		Addr <=  "00001100100100";
		Trees_din <= x"03f80604";
		wait for Clk_period;
		Addr <=  "00001100100101";
		Trees_din <= x"ffea0d65";
		wait for Clk_period;
		Addr <=  "00001100100110";
		Trees_din <= x"009a0d65";
		wait for Clk_period;
		Addr <=  "00001100100111";
		Trees_din <= x"16019d08";
		wait for Clk_period;
		Addr <=  "00001100101000";
		Trees_din <= x"05fe1904";
		wait for Clk_period;
		Addr <=  "00001100101001";
		Trees_din <= x"007a0d65";
		wait for Clk_period;
		Addr <=  "00001100101010";
		Trees_din <= x"ff960d65";
		wait for Clk_period;
		Addr <=  "00001100101011";
		Trees_din <= x"1603fe04";
		wait for Clk_period;
		Addr <=  "00001100101100";
		Trees_din <= x"00e50d65";
		wait for Clk_period;
		Addr <=  "00001100101101";
		Trees_din <= x"ffb70d65";
		wait for Clk_period;
		Addr <=  "00001100101110";
		Trees_din <= x"00167638";
		wait for Clk_period;
		Addr <=  "00001100101111";
		Trees_din <= x"03f5ed20";
		wait for Clk_period;
		Addr <=  "00001100110000";
		Trees_din <= x"0c018c10";
		wait for Clk_period;
		Addr <=  "00001100110001";
		Trees_din <= x"0b049d08";
		wait for Clk_period;
		Addr <=  "00001100110010";
		Trees_din <= x"0bf96204";
		wait for Clk_period;
		Addr <=  "00001100110011";
		Trees_din <= x"ffd70d65";
		wait for Clk_period;
		Addr <=  "00001100110100";
		Trees_din <= x"00ae0d65";
		wait for Clk_period;
		Addr <=  "00001100110101";
		Trees_din <= x"06f3f704";
		wait for Clk_period;
		Addr <=  "00001100110110";
		Trees_din <= x"ff590d65";
		wait for Clk_period;
		Addr <=  "00001100110111";
		Trees_din <= x"004a0d65";
		wait for Clk_period;
		Addr <=  "00001100111000";
		Trees_din <= x"09005a08";
		wait for Clk_period;
		Addr <=  "00001100111001";
		Trees_din <= x"09005404";
		wait for Clk_period;
		Addr <=  "00001100111010";
		Trees_din <= x"ffd00d65";
		wait for Clk_period;
		Addr <=  "00001100111011";
		Trees_din <= x"00510d65";
		wait for Clk_period;
		Addr <=  "00001100111100";
		Trees_din <= x"0d002104";
		wait for Clk_period;
		Addr <=  "00001100111101";
		Trees_din <= x"fffb0d65";
		wait for Clk_period;
		Addr <=  "00001100111110";
		Trees_din <= x"ff270d65";
		wait for Clk_period;
		Addr <=  "00001100111111";
		Trees_din <= x"0e04950c";
		wait for Clk_period;
		Addr <=  "00001101000000";
		Trees_din <= x"16040008";
		wait for Clk_period;
		Addr <=  "00001101000001";
		Trees_din <= x"17000604";
		wait for Clk_period;
		Addr <=  "00001101000010";
		Trees_din <= x"00690d65";
		wait for Clk_period;
		Addr <=  "00001101000011";
		Trees_din <= x"009f0d65";
		wait for Clk_period;
		Addr <=  "00001101000100";
		Trees_din <= x"ff9e0d65";
		wait for Clk_period;
		Addr <=  "00001101000101";
		Trees_din <= x"00148708";
		wait for Clk_period;
		Addr <=  "00001101000110";
		Trees_din <= x"0bfb1004";
		wait for Clk_period;
		Addr <=  "00001101000111";
		Trees_din <= x"00930d65";
		wait for Clk_period;
		Addr <=  "00001101001000";
		Trees_din <= x"fff10d65";
		wait for Clk_period;
		Addr <=  "00001101001001";
		Trees_din <= x"ff280d65";
		wait for Clk_period;
		Addr <=  "00001101001010";
		Trees_din <= x"010d4f0c";
		wait for Clk_period;
		Addr <=  "00001101001011";
		Trees_din <= x"0a07cb04";
		wait for Clk_period;
		Addr <=  "00001101001100";
		Trees_din <= x"00a80d65";
		wait for Clk_period;
		Addr <=  "00001101001101";
		Trees_din <= x"15009404";
		wait for Clk_period;
		Addr <=  "00001101001110";
		Trees_din <= x"ffc30d65";
		wait for Clk_period;
		Addr <=  "00001101001111";
		Trees_din <= x"007e0d65";
		wait for Clk_period;
		Addr <=  "00001101010000";
		Trees_din <= x"0bf88604";
		wait for Clk_period;
		Addr <=  "00001101010001";
		Trees_din <= x"ffa70d65";
		wait for Clk_period;
		Addr <=  "00001101010010";
		Trees_din <= x"07005508";
		wait for Clk_period;
		Addr <=  "00001101010011";
		Trees_din <= x"1a00db04";
		wait for Clk_period;
		Addr <=  "00001101010100";
		Trees_din <= x"ffd30d65";
		wait for Clk_period;
		Addr <=  "00001101010101";
		Trees_din <= x"00910d65";
		wait for Clk_period;
		Addr <=  "00001101010110";
		Trees_din <= x"020a7304";
		wait for Clk_period;
		Addr <=  "00001101010111";
		Trees_din <= x"00a20d65";
		wait for Clk_period;
		Addr <=  "00001101011000";
		Trees_din <= x"fffc0d65";
		wait for Clk_period;
		Addr <=  "00001101011001";
		Trees_din <= x"00119250";
		wait for Clk_period;
		Addr <=  "00001101011010";
		Trees_din <= x"0003aa2c";
		wait for Clk_period;
		Addr <=  "00001101011011";
		Trees_din <= x"01fdfc18";
		wait for Clk_period;
		Addr <=  "00001101011100";
		Trees_din <= x"0c01ef10";
		wait for Clk_period;
		Addr <=  "00001101011101";
		Trees_din <= x"00015508";
		wait for Clk_period;
		Addr <=  "00001101011110";
		Trees_din <= x"05fdb604";
		wait for Clk_period;
		Addr <=  "00001101011111";
		Trees_din <= x"ff730eb1";
		wait for Clk_period;
		Addr <=  "00001101100000";
		Trees_din <= x"00630eb1";
		wait for Clk_period;
		Addr <=  "00001101100001";
		Trees_din <= x"06f69704";
		wait for Clk_period;
		Addr <=  "00001101100010";
		Trees_din <= x"016a0eb1";
		wait for Clk_period;
		Addr <=  "00001101100011";
		Trees_din <= x"00110eb1";
		wait for Clk_period;
		Addr <=  "00001101100100";
		Trees_din <= x"1900b004";
		wait for Clk_period;
		Addr <=  "00001101100101";
		Trees_din <= x"ff6d0eb1";
		wait for Clk_period;
		Addr <=  "00001101100110";
		Trees_din <= x"001e0eb1";
		wait for Clk_period;
		Addr <=  "00001101100111";
		Trees_din <= x"1b006610";
		wait for Clk_period;
		Addr <=  "00001101101000";
		Trees_din <= x"0bf98508";
		wait for Clk_period;
		Addr <=  "00001101101001";
		Trees_din <= x"12023f04";
		wait for Clk_period;
		Addr <=  "00001101101010";
		Trees_din <= x"ff760eb1";
		wait for Clk_period;
		Addr <=  "00001101101011";
		Trees_din <= x"00ac0eb1";
		wait for Clk_period;
		Addr <=  "00001101101100";
		Trees_din <= x"1603fe04";
		wait for Clk_period;
		Addr <=  "00001101101101";
		Trees_din <= x"ff760eb1";
		wait for Clk_period;
		Addr <=  "00001101101110";
		Trees_din <= x"00170eb1";
		wait for Clk_period;
		Addr <=  "00001101101111";
		Trees_din <= x"00770eb1";
		wait for Clk_period;
		Addr <=  "00001101110000";
		Trees_din <= x"02107e1c";
		wait for Clk_period;
		Addr <=  "00001101110001";
		Trees_din <= x"0113e910";
		wait for Clk_period;
		Addr <=  "00001101110010";
		Trees_din <= x"09005d08";
		wait for Clk_period;
		Addr <=  "00001101110011";
		Trees_din <= x"0007fa04";
		wait for Clk_period;
		Addr <=  "00001101110100";
		Trees_din <= x"fffa0eb1";
		wait for Clk_period;
		Addr <=  "00001101110101";
		Trees_din <= x"00350eb1";
		wait for Clk_period;
		Addr <=  "00001101110110";
		Trees_din <= x"0d00ef04";
		wait for Clk_period;
		Addr <=  "00001101110111";
		Trees_din <= x"01310eb1";
		wait for Clk_period;
		Addr <=  "00001101111000";
		Trees_din <= x"00510eb1";
		wait for Clk_period;
		Addr <=  "00001101111001";
		Trees_din <= x"0efa8a08";
		wait for Clk_period;
		Addr <=  "00001101111010";
		Trees_din <= x"000e4f04";
		wait for Clk_period;
		Addr <=  "00001101111011";
		Trees_din <= x"ffad0eb1";
		wait for Clk_period;
		Addr <=  "00001101111100";
		Trees_din <= x"00bd0eb1";
		wait for Clk_period;
		Addr <=  "00001101111101";
		Trees_din <= x"ff6e0eb1";
		wait for Clk_period;
		Addr <=  "00001101111110";
		Trees_din <= x"06f68504";
		wait for Clk_period;
		Addr <=  "00001101111111";
		Trees_din <= x"ff6e0eb1";
		wait for Clk_period;
		Addr <=  "00001110000000";
		Trees_din <= x"003b0eb1";
		wait for Clk_period;
		Addr <=  "00001110000001";
		Trees_din <= x"00167638";
		wait for Clk_period;
		Addr <=  "00001110000010";
		Trees_din <= x"03f6251c";
		wait for Clk_period;
		Addr <=  "00001110000011";
		Trees_din <= x"0c018c10";
		wait for Clk_period;
		Addr <=  "00001110000100";
		Trees_din <= x"0f000708";
		wait for Clk_period;
		Addr <=  "00001110000101";
		Trees_din <= x"19007704";
		wait for Clk_period;
		Addr <=  "00001110000110";
		Trees_din <= x"00850eb1";
		wait for Clk_period;
		Addr <=  "00001110000111";
		Trees_din <= x"ff8f0eb1";
		wait for Clk_period;
		Addr <=  "00001110001000";
		Trees_din <= x"0b049d04";
		wait for Clk_period;
		Addr <=  "00001110001001";
		Trees_din <= x"009f0eb1";
		wait for Clk_period;
		Addr <=  "00001110001010";
		Trees_din <= x"00180eb1";
		wait for Clk_period;
		Addr <=  "00001110001011";
		Trees_din <= x"04faf608";
		wait for Clk_period;
		Addr <=  "00001110001100";
		Trees_din <= x"04f93f04";
		wait for Clk_period;
		Addr <=  "00001110001101";
		Trees_din <= x"001b0eb1";
		wait for Clk_period;
		Addr <=  "00001110001110";
		Trees_din <= x"ff7e0eb1";
		wait for Clk_period;
		Addr <=  "00001110001111";
		Trees_din <= x"00a00eb1";
		wait for Clk_period;
		Addr <=  "00001110010000";
		Trees_din <= x"1700060c";
		wait for Clk_period;
		Addr <=  "00001110010001";
		Trees_din <= x"11009a04";
		wait for Clk_period;
		Addr <=  "00001110010010";
		Trees_din <= x"00ab0eb1";
		wait for Clk_period;
		Addr <=  "00001110010011";
		Trees_din <= x"0f000004";
		wait for Clk_period;
		Addr <=  "00001110010100";
		Trees_din <= x"ff4e0eb1";
		wait for Clk_period;
		Addr <=  "00001110010101";
		Trees_din <= x"003f0eb1";
		wait for Clk_period;
		Addr <=  "00001110010110";
		Trees_din <= x"0a036d08";
		wait for Clk_period;
		Addr <=  "00001110010111";
		Trees_din <= x"04f55a04";
		wait for Clk_period;
		Addr <=  "00001110011000";
		Trees_din <= x"000d0eb1";
		wait for Clk_period;
		Addr <=  "00001110011001";
		Trees_din <= x"00a10eb1";
		wait for Clk_period;
		Addr <=  "00001110011010";
		Trees_din <= x"09004c04";
		wait for Clk_period;
		Addr <=  "00001110011011";
		Trees_din <= x"ff480eb1";
		wait for Clk_period;
		Addr <=  "00001110011100";
		Trees_din <= x"00600eb1";
		wait for Clk_period;
		Addr <=  "00001110011101";
		Trees_din <= x"010d4f0c";
		wait for Clk_period;
		Addr <=  "00001110011110";
		Trees_din <= x"0a07cb04";
		wait for Clk_period;
		Addr <=  "00001110011111";
		Trees_din <= x"00a40eb1";
		wait for Clk_period;
		Addr <=  "00001110100000";
		Trees_din <= x"02028904";
		wait for Clk_period;
		Addr <=  "00001110100001";
		Trees_din <= x"00740eb1";
		wait for Clk_period;
		Addr <=  "00001110100010";
		Trees_din <= x"ffc30eb1";
		wait for Clk_period;
		Addr <=  "00001110100011";
		Trees_din <= x"0bf88604";
		wait for Clk_period;
		Addr <=  "00001110100100";
		Trees_din <= x"ffa70eb1";
		wait for Clk_period;
		Addr <=  "00001110100101";
		Trees_din <= x"07005508";
		wait for Clk_period;
		Addr <=  "00001110100110";
		Trees_din <= x"1a00db04";
		wait for Clk_period;
		Addr <=  "00001110100111";
		Trees_din <= x"ffd10eb1";
		wait for Clk_period;
		Addr <=  "00001110101000";
		Trees_din <= x"00860eb1";
		wait for Clk_period;
		Addr <=  "00001110101001";
		Trees_din <= x"1f000204";
		wait for Clk_period;
		Addr <=  "00001110101010";
		Trees_din <= x"009a0eb1";
		wait for Clk_period;
		Addr <=  "00001110101011";
		Trees_din <= x"ffef0eb1";
		wait for Clk_period;
		Addr <=  "00001110101100";
		Trees_din <= x"00153268";
		wait for Clk_period;
		Addr <=  "00001110101101";
		Trees_din <= x"00058428";
		wait for Clk_period;
		Addr <=  "00001110101110";
		Trees_din <= x"1f000014";
		wait for Clk_period;
		Addr <=  "00001110101111";
		Trees_din <= x"00fe7b04";
		wait for Clk_period;
		Addr <=  "00001110110000";
		Trees_din <= x"ff69100d";
		wait for Clk_period;
		Addr <=  "00001110110001";
		Trees_din <= x"01fd7808";
		wait for Clk_period;
		Addr <=  "00001110110010";
		Trees_din <= x"07005804";
		wait for Clk_period;
		Addr <=  "00001110110011";
		Trees_din <= x"0072100d";
		wait for Clk_period;
		Addr <=  "00001110110100";
		Trees_din <= x"ff92100d";
		wait for Clk_period;
		Addr <=  "00001110110101";
		Trees_din <= x"04060d04";
		wait for Clk_period;
		Addr <=  "00001110110110";
		Trees_din <= x"ff9b100d";
		wait for Clk_period;
		Addr <=  "00001110110111";
		Trees_din <= x"0002100d";
		wait for Clk_period;
		Addr <=  "00001110111000";
		Trees_din <= x"0f005810";
		wait for Clk_period;
		Addr <=  "00001110111001";
		Trees_din <= x"09005008";
		wait for Clk_period;
		Addr <=  "00001110111010";
		Trees_din <= x"13014d04";
		wait for Clk_period;
		Addr <=  "00001110111011";
		Trees_din <= x"ff8a100d";
		wait for Clk_period;
		Addr <=  "00001110111100";
		Trees_din <= x"001f100d";
		wait for Clk_period;
		Addr <=  "00001110111101";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00001110111110";
		Trees_din <= x"0184100d";
		wait for Clk_period;
		Addr <=  "00001110111111";
		Trees_din <= x"004c100d";
		wait for Clk_period;
		Addr <=  "00001111000000";
		Trees_din <= x"ff79100d";
		wait for Clk_period;
		Addr <=  "00001111000001";
		Trees_din <= x"0101df20";
		wait for Clk_period;
		Addr <=  "00001111000010";
		Trees_din <= x"05005810";
		wait for Clk_period;
		Addr <=  "00001111000011";
		Trees_din <= x"13f8dd08";
		wait for Clk_period;
		Addr <=  "00001111000100";
		Trees_din <= x"16014004";
		wait for Clk_period;
		Addr <=  "00001111000101";
		Trees_din <= x"ff36100d";
		wait for Clk_period;
		Addr <=  "00001111000110";
		Trees_din <= x"003c100d";
		wait for Clk_period;
		Addr <=  "00001111000111";
		Trees_din <= x"10fa9004";
		wait for Clk_period;
		Addr <=  "00001111001000";
		Trees_din <= x"0028100d";
		wait for Clk_period;
		Addr <=  "00001111001001";
		Trees_din <= x"0091100d";
		wait for Clk_period;
		Addr <=  "00001111001010";
		Trees_din <= x"00103308";
		wait for Clk_period;
		Addr <=  "00001111001011";
		Trees_din <= x"11044a04";
		wait for Clk_period;
		Addr <=  "00001111001100";
		Trees_din <= x"ff96100d";
		wait for Clk_period;
		Addr <=  "00001111001101";
		Trees_din <= x"008a100d";
		wait for Clk_period;
		Addr <=  "00001111001110";
		Trees_din <= x"15008104";
		wait for Clk_period;
		Addr <=  "00001111001111";
		Trees_din <= x"ffa8100d";
		wait for Clk_period;
		Addr <=  "00001111010000";
		Trees_din <= x"0098100d";
		wait for Clk_period;
		Addr <=  "00001111010001";
		Trees_din <= x"06f34c10";
		wait for Clk_period;
		Addr <=  "00001111010010";
		Trees_din <= x"0203d008";
		wait for Clk_period;
		Addr <=  "00001111010011";
		Trees_din <= x"07005c04";
		wait for Clk_period;
		Addr <=  "00001111010100";
		Trees_din <= x"00be100d";
		wait for Clk_period;
		Addr <=  "00001111010101";
		Trees_din <= x"ffda100d";
		wait for Clk_period;
		Addr <=  "00001111010110";
		Trees_din <= x"0afd6404";
		wait for Clk_period;
		Addr <=  "00001111010111";
		Trees_din <= x"ffe8100d";
		wait for Clk_period;
		Addr <=  "00001111011000";
		Trees_din <= x"0074100d";
		wait for Clk_period;
		Addr <=  "00001111011001";
		Trees_din <= x"000b5608";
		wait for Clk_period;
		Addr <=  "00001111011010";
		Trees_din <= x"1003c104";
		wait for Clk_period;
		Addr <=  "00001111011011";
		Trees_din <= x"0015100d";
		wait for Clk_period;
		Addr <=  "00001111011100";
		Trees_din <= x"ffa0100d";
		wait for Clk_period;
		Addr <=  "00001111011101";
		Trees_din <= x"010a1f04";
		wait for Clk_period;
		Addr <=  "00001111011110";
		Trees_din <= x"004d100d";
		wait for Clk_period;
		Addr <=  "00001111011111";
		Trees_din <= x"000a100d";
		wait for Clk_period;
		Addr <=  "00001111100000";
		Trees_din <= x"010d4f1c";
		wait for Clk_period;
		Addr <=  "00001111100001";
		Trees_din <= x"020d0614";
		wait for Clk_period;
		Addr <=  "00001111100010";
		Trees_din <= x"1a013710";
		wait for Clk_period;
		Addr <=  "00001111100011";
		Trees_din <= x"0a07cb08";
		wait for Clk_period;
		Addr <=  "00001111100100";
		Trees_din <= x"03faba04";
		wait for Clk_period;
		Addr <=  "00001111100101";
		Trees_din <= x"009f100d";
		wait for Clk_period;
		Addr <=  "00001111100110";
		Trees_din <= x"004f100d";
		wait for Clk_period;
		Addr <=  "00001111100111";
		Trees_din <= x"1c003104";
		wait for Clk_period;
		Addr <=  "00001111101000";
		Trees_din <= x"ffc8100d";
		wait for Clk_period;
		Addr <=  "00001111101001";
		Trees_din <= x"006c100d";
		wait for Clk_period;
		Addr <=  "00001111101010";
		Trees_din <= x"000e100d";
		wait for Clk_period;
		Addr <=  "00001111101011";
		Trees_din <= x"03f26104";
		wait for Clk_period;
		Addr <=  "00001111101100";
		Trees_din <= x"001b100d";
		wait for Clk_period;
		Addr <=  "00001111101101";
		Trees_din <= x"fff1100d";
		wait for Clk_period;
		Addr <=  "00001111101110";
		Trees_din <= x"00192f18";
		wait for Clk_period;
		Addr <=  "00001111101111";
		Trees_din <= x"03f2890c";
		wait for Clk_period;
		Addr <=  "00001111110000";
		Trees_din <= x"06f3a804";
		wait for Clk_period;
		Addr <=  "00001111110001";
		Trees_din <= x"006e100d";
		wait for Clk_period;
		Addr <=  "00001111110010";
		Trees_din <= x"12028804";
		wait for Clk_period;
		Addr <=  "00001111110011";
		Trees_din <= x"ff3b100d";
		wait for Clk_period;
		Addr <=  "00001111110100";
		Trees_din <= x"0029100d";
		wait for Clk_period;
		Addr <=  "00001111110101";
		Trees_din <= x"0c03d208";
		wait for Clk_period;
		Addr <=  "00001111110110";
		Trees_din <= x"1a00d704";
		wait for Clk_period;
		Addr <=  "00001111110111";
		Trees_din <= x"008d100d";
		wait for Clk_period;
		Addr <=  "00001111111000";
		Trees_din <= x"fffb100d";
		wait for Clk_period;
		Addr <=  "00001111111001";
		Trees_din <= x"ff5d100d";
		wait for Clk_period;
		Addr <=  "00001111111010";
		Trees_din <= x"03f4e80c";
		wait for Clk_period;
		Addr <=  "00001111111011";
		Trees_din <= x"19008908";
		wait for Clk_period;
		Addr <=  "00001111111100";
		Trees_din <= x"09004f04";
		wait for Clk_period;
		Addr <=  "00001111111101";
		Trees_din <= x"ff44100d";
		wait for Clk_period;
		Addr <=  "00001111111110";
		Trees_din <= x"008a100d";
		wait for Clk_period;
		Addr <=  "00001111111111";
		Trees_din <= x"009c100d";
		wait for Clk_period;
		Addr <=  "00010000000000";
		Trees_din <= x"001b5104";
		wait for Clk_period;
		Addr <=  "00010000000001";
		Trees_din <= x"005e100d";
		wait for Clk_period;
		Addr <=  "00010000000010";
		Trees_din <= x"ff70100d";
		wait for Clk_period;
		Addr <=  "00010000000011";
		Trees_din <= x"00167668";
		wait for Clk_period;
		Addr <=  "00010000000100";
		Trees_din <= x"0003aa2c";
		wait for Clk_period;
		Addr <=  "00010000000101";
		Trees_din <= x"01fdfc18";
		wait for Clk_period;
		Addr <=  "00010000000110";
		Trees_din <= x"0c01ef10";
		wait for Clk_period;
		Addr <=  "00010000000111";
		Trees_din <= x"0c014408";
		wait for Clk_period;
		Addr <=  "00010000001000";
		Trees_din <= x"0c007c04";
		wait for Clk_period;
		Addr <=  "00010000001001";
		Trees_din <= x"00361149";
		wait for Clk_period;
		Addr <=  "00010000001010";
		Trees_din <= x"ff771149";
		wait for Clk_period;
		Addr <=  "00010000001011";
		Trees_din <= x"12010604";
		wait for Clk_period;
		Addr <=  "00010000001100";
		Trees_din <= x"ff9d1149";
		wait for Clk_period;
		Addr <=  "00010000001101";
		Trees_din <= x"01041149";
		wait for Clk_period;
		Addr <=  "00010000001110";
		Trees_din <= x"0408ca04";
		wait for Clk_period;
		Addr <=  "00010000001111";
		Trees_din <= x"ff721149";
		wait for Clk_period;
		Addr <=  "00010000010000";
		Trees_din <= x"00291149";
		wait for Clk_period;
		Addr <=  "00010000010001";
		Trees_din <= x"1b006610";
		wait for Clk_period;
		Addr <=  "00010000010010";
		Trees_din <= x"08022008";
		wait for Clk_period;
		Addr <=  "00010000010011";
		Trees_din <= x"1e009504";
		wait for Clk_period;
		Addr <=  "00010000010100";
		Trees_din <= x"ff771149";
		wait for Clk_period;
		Addr <=  "00010000010101";
		Trees_din <= x"00351149";
		wait for Clk_period;
		Addr <=  "00010000010110";
		Trees_din <= x"08024004";
		wait for Clk_period;
		Addr <=  "00010000010111";
		Trees_din <= x"00d81149";
		wait for Clk_period;
		Addr <=  "00010000011000";
		Trees_din <= x"ff901149";
		wait for Clk_period;
		Addr <=  "00010000011001";
		Trees_din <= x"00711149";
		wait for Clk_period;
		Addr <=  "00010000011010";
		Trees_din <= x"000f6f1c";
		wait for Clk_period;
		Addr <=  "00010000011011";
		Trees_din <= x"09005d10";
		wait for Clk_period;
		Addr <=  "00010000011100";
		Trees_din <= x"06f76d08";
		wait for Clk_period;
		Addr <=  "00010000011101";
		Trees_din <= x"02ff5104";
		wait for Clk_period;
		Addr <=  "00010000011110";
		Trees_din <= x"00831149";
		wait for Clk_period;
		Addr <=  "00010000011111";
		Trees_din <= x"00141149";
		wait for Clk_period;
		Addr <=  "00010000100000";
		Trees_din <= x"01029904";
		wait for Clk_period;
		Addr <=  "00010000100001";
		Trees_din <= x"00221149";
		wait for Clk_period;
		Addr <=  "00010000100010";
		Trees_din <= x"ffc21149";
		wait for Clk_period;
		Addr <=  "00010000100011";
		Trees_din <= x"09005f08";
		wait for Clk_period;
		Addr <=  "00010000100100";
		Trees_din <= x"04ffda04";
		wait for Clk_period;
		Addr <=  "00010000100101";
		Trees_din <= x"00fb1149";
		wait for Clk_period;
		Addr <=  "00010000100110";
		Trees_din <= x"00161149";
		wait for Clk_period;
		Addr <=  "00010000100111";
		Trees_din <= x"ffcd1149";
		wait for Clk_period;
		Addr <=  "00010000101000";
		Trees_din <= x"0c033110";
		wait for Clk_period;
		Addr <=  "00010000101001";
		Trees_din <= x"0205a108";
		wait for Clk_period;
		Addr <=  "00010000101010";
		Trees_din <= x"1703f804";
		wait for Clk_period;
		Addr <=  "00010000101011";
		Trees_din <= x"00671149";
		wait for Clk_period;
		Addr <=  "00010000101100";
		Trees_din <= x"ffb91149";
		wait for Clk_period;
		Addr <=  "00010000101101";
		Trees_din <= x"16039c04";
		wait for Clk_period;
		Addr <=  "00010000101110";
		Trees_din <= x"ffef1149";
		wait for Clk_period;
		Addr <=  "00010000101111";
		Trees_din <= x"00681149";
		wait for Clk_period;
		Addr <=  "00010000110000";
		Trees_din <= x"1e007808";
		wait for Clk_period;
		Addr <=  "00010000110001";
		Trees_din <= x"18003b04";
		wait for Clk_period;
		Addr <=  "00010000110010";
		Trees_din <= x"00831149";
		wait for Clk_period;
		Addr <=  "00010000110011";
		Trees_din <= x"ffb81149";
		wait for Clk_period;
		Addr <=  "00010000110100";
		Trees_din <= x"0f000004";
		wait for Clk_period;
		Addr <=  "00010000110101";
		Trees_din <= x"ff5d1149";
		wait for Clk_period;
		Addr <=  "00010000110110";
		Trees_din <= x"00951149";
		wait for Clk_period;
		Addr <=  "00010000110111";
		Trees_din <= x"010d4f14";
		wait for Clk_period;
		Addr <=  "00010000111000";
		Trees_din <= x"0a07cb0c";
		wait for Clk_period;
		Addr <=  "00010000111001";
		Trees_din <= x"0d000008";
		wait for Clk_period;
		Addr <=  "00010000111010";
		Trees_din <= x"18003e04";
		wait for Clk_period;
		Addr <=  "00010000111011";
		Trees_din <= x"ffc11149";
		wait for Clk_period;
		Addr <=  "00010000111100";
		Trees_din <= x"00821149";
		wait for Clk_period;
		Addr <=  "00010000111101";
		Trees_din <= x"009e1149";
		wait for Clk_period;
		Addr <=  "00010000111110";
		Trees_din <= x"1a00df04";
		wait for Clk_period;
		Addr <=  "00010000111111";
		Trees_din <= x"00621149";
		wait for Clk_period;
		Addr <=  "00010001000000";
		Trees_din <= x"ffc21149";
		wait for Clk_period;
		Addr <=  "00010001000001";
		Trees_din <= x"0bf88604";
		wait for Clk_period;
		Addr <=  "00010001000010";
		Trees_din <= x"ffa11149";
		wait for Clk_period;
		Addr <=  "00010001000011";
		Trees_din <= x"07005510";
		wait for Clk_period;
		Addr <=  "00010001000100";
		Trees_din <= x"1a00db08";
		wait for Clk_period;
		Addr <=  "00010001000101";
		Trees_din <= x"1c004004";
		wait for Clk_period;
		Addr <=  "00010001000110";
		Trees_din <= x"ff741149";
		wait for Clk_period;
		Addr <=  "00010001000111";
		Trees_din <= x"00731149";
		wait for Clk_period;
		Addr <=  "00010001001000";
		Trees_din <= x"0018ac04";
		wait for Clk_period;
		Addr <=  "00010001001001";
		Trees_din <= x"00191149";
		wait for Clk_period;
		Addr <=  "00010001001010";
		Trees_din <= x"008a1149";
		wait for Clk_period;
		Addr <=  "00010001001011";
		Trees_din <= x"020a7308";
		wait for Clk_period;
		Addr <=  "00010001001100";
		Trees_din <= x"01164204";
		wait for Clk_period;
		Addr <=  "00010001001101";
		Trees_din <= x"009d1149";
		wait for Clk_period;
		Addr <=  "00010001001110";
		Trees_din <= x"ffe51149";
		wait for Clk_period;
		Addr <=  "00010001001111";
		Trees_din <= x"17000804";
		wait for Clk_period;
		Addr <=  "00010001010000";
		Trees_din <= x"00541149";
		wait for Clk_period;
		Addr <=  "00010001010001";
		Trees_din <= x"ff6a1149";
		wait for Clk_period;
		Addr <=  "00010001010010";
		Trees_din <= x"00167674";
		wait for Clk_period;
		Addr <=  "00010001010011";
		Trees_din <= x"0007903c";
		wait for Clk_period;
		Addr <=  "00010001010100";
		Trees_din <= x"0000af1c";
		wait for Clk_period;
		Addr <=  "00010001010101";
		Trees_din <= x"02fba50c";
		wait for Clk_period;
		Addr <=  "00010001010110";
		Trees_din <= x"14003304";
		wait for Clk_period;
		Addr <=  "00010001010111";
		Trees_din <= x"00b612a5";
		wait for Clk_period;
		Addr <=  "00010001011000";
		Trees_din <= x"1e005e04";
		wait for Clk_period;
		Addr <=  "00010001011001";
		Trees_din <= x"001212a5";
		wait for Clk_period;
		Addr <=  "00010001011010";
		Trees_din <= x"ffa412a5";
		wait for Clk_period;
		Addr <=  "00010001011011";
		Trees_din <= x"10f8a608";
		wait for Clk_period;
		Addr <=  "00010001011100";
		Trees_din <= x"1a00cc04";
		wait for Clk_period;
		Addr <=  "00010001011101";
		Trees_din <= x"00d512a5";
		wait for Clk_period;
		Addr <=  "00010001011110";
		Trees_din <= x"ff9c12a5";
		wait for Clk_period;
		Addr <=  "00010001011111";
		Trees_din <= x"1e004a04";
		wait for Clk_period;
		Addr <=  "00010001100000";
		Trees_din <= x"004912a5";
		wait for Clk_period;
		Addr <=  "00010001100001";
		Trees_din <= x"ff6912a5";
		wait for Clk_period;
		Addr <=  "00010001100010";
		Trees_din <= x"03fe2510";
		wait for Clk_period;
		Addr <=  "00010001100011";
		Trees_din <= x"13ffcc08";
		wait for Clk_period;
		Addr <=  "00010001100100";
		Trees_din <= x"13f8dd04";
		wait for Clk_period;
		Addr <=  "00010001100101";
		Trees_din <= x"003112a5";
		wait for Clk_period;
		Addr <=  "00010001100110";
		Trees_din <= x"ff7312a5";
		wait for Clk_period;
		Addr <=  "00010001100111";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00010001101000";
		Trees_din <= x"00b312a5";
		wait for Clk_period;
		Addr <=  "00010001101001";
		Trees_din <= x"ffb412a5";
		wait for Clk_period;
		Addr <=  "00010001101010";
		Trees_din <= x"1201f608";
		wait for Clk_period;
		Addr <=  "00010001101011";
		Trees_din <= x"0e021e04";
		wait for Clk_period;
		Addr <=  "00010001101100";
		Trees_din <= x"ffc712a5";
		wait for Clk_period;
		Addr <=  "00010001101101";
		Trees_din <= x"005b12a5";
		wait for Clk_period;
		Addr <=  "00010001101110";
		Trees_din <= x"1b004004";
		wait for Clk_period;
		Addr <=  "00010001101111";
		Trees_din <= x"000812a5";
		wait for Clk_period;
		Addr <=  "00010001110000";
		Trees_din <= x"00a212a5";
		wait for Clk_period;
		Addr <=  "00010001110001";
		Trees_din <= x"04ff5720";
		wait for Clk_period;
		Addr <=  "00010001110010";
		Trees_din <= x"00119210";
		wait for Clk_period;
		Addr <=  "00010001110011";
		Trees_din <= x"01037508";
		wait for Clk_period;
		Addr <=  "00010001110100";
		Trees_din <= x"05fff704";
		wait for Clk_period;
		Addr <=  "00010001110101";
		Trees_din <= x"006312a5";
		wait for Clk_period;
		Addr <=  "00010001110110";
		Trees_din <= x"ffd512a5";
		wait for Clk_period;
		Addr <=  "00010001110111";
		Trees_din <= x"0afd4004";
		wait for Clk_period;
		Addr <=  "00010001111000";
		Trees_din <= x"ffda12a5";
		wait for Clk_period;
		Addr <=  "00010001111001";
		Trees_din <= x"002012a5";
		wait for Clk_period;
		Addr <=  "00010001111010";
		Trees_din <= x"0c028808";
		wait for Clk_period;
		Addr <=  "00010001111011";
		Trees_din <= x"0203d004";
		wait for Clk_period;
		Addr <=  "00010001111100";
		Trees_din <= x"007c12a5";
		wait for Clk_period;
		Addr <=  "00010001111101";
		Trees_din <= x"002a12a5";
		wait for Clk_period;
		Addr <=  "00010001111110";
		Trees_din <= x"1b003a04";
		wait for Clk_period;
		Addr <=  "00010001111111";
		Trees_din <= x"ffd612a5";
		wait for Clk_period;
		Addr <=  "00010010000000";
		Trees_din <= x"004912a5";
		wait for Clk_period;
		Addr <=  "00010010000001";
		Trees_din <= x"1c004d10";
		wait for Clk_period;
		Addr <=  "00010010000010";
		Trees_din <= x"18003d08";
		wait for Clk_period;
		Addr <=  "00010010000011";
		Trees_din <= x"0e002f04";
		wait for Clk_period;
		Addr <=  "00010010000100";
		Trees_din <= x"ffb712a5";
		wait for Clk_period;
		Addr <=  "00010010000101";
		Trees_din <= x"005d12a5";
		wait for Clk_period;
		Addr <=  "00010010000110";
		Trees_din <= x"0afb1504";
		wait for Clk_period;
		Addr <=  "00010010000111";
		Trees_din <= x"000812a5";
		wait for Clk_period;
		Addr <=  "00010010001000";
		Trees_din <= x"00b012a5";
		wait for Clk_period;
		Addr <=  "00010010001001";
		Trees_din <= x"01042f04";
		wait for Clk_period;
		Addr <=  "00010010001010";
		Trees_din <= x"000b12a5";
		wait for Clk_period;
		Addr <=  "00010010001011";
		Trees_din <= x"ff3e12a5";
		wait for Clk_period;
		Addr <=  "00010010001100";
		Trees_din <= x"010d4f1c";
		wait for Clk_period;
		Addr <=  "00010010001101";
		Trees_din <= x"0a07cb14";
		wait for Clk_period;
		Addr <=  "00010010001110";
		Trees_din <= x"0d000008";
		wait for Clk_period;
		Addr <=  "00010010001111";
		Trees_din <= x"05fd8604";
		wait for Clk_period;
		Addr <=  "00010010010000";
		Trees_din <= x"007b12a5";
		wait for Clk_period;
		Addr <=  "00010010010001";
		Trees_din <= x"ffbb12a5";
		wait for Clk_period;
		Addr <=  "00010010010010";
		Trees_din <= x"1f000c04";
		wait for Clk_period;
		Addr <=  "00010010010011";
		Trees_din <= x"009c12a5";
		wait for Clk_period;
		Addr <=  "00010010010100";
		Trees_din <= x"03f06b04";
		wait for Clk_period;
		Addr <=  "00010010010101";
		Trees_din <= x"ffb712a5";
		wait for Clk_period;
		Addr <=  "00010010010110";
		Trees_din <= x"008212a5";
		wait for Clk_period;
		Addr <=  "00010010010111";
		Trees_din <= x"08015704";
		wait for Clk_period;
		Addr <=  "00010010011000";
		Trees_din <= x"ffc412a5";
		wait for Clk_period;
		Addr <=  "00010010011001";
		Trees_din <= x"005b12a5";
		wait for Clk_period;
		Addr <=  "00010010011010";
		Trees_din <= x"001be914";
		wait for Clk_period;
		Addr <=  "00010010011011";
		Trees_din <= x"0bf95b08";
		wait for Clk_period;
		Addr <=  "00010010011100";
		Trees_din <= x"18003d04";
		wait for Clk_period;
		Addr <=  "00010010011101";
		Trees_din <= x"ff3b12a5";
		wait for Clk_period;
		Addr <=  "00010010011110";
		Trees_din <= x"ffd412a5";
		wait for Clk_period;
		Addr <=  "00010010011111";
		Trees_din <= x"03f7b308";
		wait for Clk_period;
		Addr <=  "00010010100000";
		Trees_din <= x"03f09e04";
		wait for Clk_period;
		Addr <=  "00010010100001";
		Trees_din <= x"ff9712a5";
		wait for Clk_period;
		Addr <=  "00010010100010";
		Trees_din <= x"006212a5";
		wait for Clk_period;
		Addr <=  "00010010100011";
		Trees_din <= x"ff9b12a5";
		wait for Clk_period;
		Addr <=  "00010010100100";
		Trees_din <= x"1302d208";
		wait for Clk_period;
		Addr <=  "00010010100101";
		Trees_din <= x"0802cf04";
		wait for Clk_period;
		Addr <=  "00010010100110";
		Trees_din <= x"009612a5";
		wait for Clk_period;
		Addr <=  "00010010100111";
		Trees_din <= x"002112a5";
		wait for Clk_period;
		Addr <=  "00010010101000";
		Trees_din <= x"ffe412a5";
		wait for Clk_period;
		Addr <=  "00010010101001";
		Trees_din <= x"0016766c";
		wait for Clk_period;
		Addr <=  "00010010101010";
		Trees_din <= x"0003aa2c";
		wait for Clk_period;
		Addr <=  "00010010101011";
		Trees_din <= x"1b003d18";
		wait for Clk_period;
		Addr <=  "00010010101100";
		Trees_din <= x"1f00000c";
		wait for Clk_period;
		Addr <=  "00010010101101";
		Trees_din <= x"0bf8e904";
		wait for Clk_period;
		Addr <=  "00010010101110";
		Trees_din <= x"003913f9";
		wait for Clk_period;
		Addr <=  "00010010101111";
		Trees_din <= x"10f72e04";
		wait for Clk_period;
		Addr <=  "00010010110000";
		Trees_din <= x"001813f9";
		wait for Clk_period;
		Addr <=  "00010010110001";
		Trees_din <= x"ff7213f9";
		wait for Clk_period;
		Addr <=  "00010010110010";
		Trees_din <= x"1f000208";
		wait for Clk_period;
		Addr <=  "00010010110011";
		Trees_din <= x"0e00c804";
		wait for Clk_period;
		Addr <=  "00010010110100";
		Trees_din <= x"ffa413f9";
		wait for Clk_period;
		Addr <=  "00010010110101";
		Trees_din <= x"00b613f9";
		wait for Clk_period;
		Addr <=  "00010010110110";
		Trees_din <= x"ff8f13f9";
		wait for Clk_period;
		Addr <=  "00010010110111";
		Trees_din <= x"0700580c";
		wait for Clk_period;
		Addr <=  "00010010111000";
		Trees_din <= x"00fe7b04";
		wait for Clk_period;
		Addr <=  "00010010111001";
		Trees_din <= x"ff8f13f9";
		wait for Clk_period;
		Addr <=  "00010010111010";
		Trees_din <= x"08001a04";
		wait for Clk_period;
		Addr <=  "00010010111011";
		Trees_din <= x"ff9413f9";
		wait for Clk_period;
		Addr <=  "00010010111100";
		Trees_din <= x"00a213f9";
		wait for Clk_period;
		Addr <=  "00010010111101";
		Trees_din <= x"09003c04";
		wait for Clk_period;
		Addr <=  "00010010111110";
		Trees_din <= x"005513f9";
		wait for Clk_period;
		Addr <=  "00010010111111";
		Trees_din <= x"ff7213f9";
		wait for Clk_period;
		Addr <=  "00010011000000";
		Trees_din <= x"1900a620";
		wait for Clk_period;
		Addr <=  "00010011000001";
		Trees_din <= x"1b003410";
		wait for Clk_period;
		Addr <=  "00010011000010";
		Trees_din <= x"11043808";
		wait for Clk_period;
		Addr <=  "00010011000011";
		Trees_din <= x"00054504";
		wait for Clk_period;
		Addr <=  "00010011000100";
		Trees_din <= x"00d513f9";
		wait for Clk_period;
		Addr <=  "00010011000101";
		Trees_din <= x"ffec13f9";
		wait for Clk_period;
		Addr <=  "00010011000110";
		Trees_din <= x"1e005f04";
		wait for Clk_period;
		Addr <=  "00010011000111";
		Trees_din <= x"ff0113f9";
		wait for Clk_period;
		Addr <=  "00010011001000";
		Trees_din <= x"003213f9";
		wait for Clk_period;
		Addr <=  "00010011001001";
		Trees_din <= x"11047908";
		wait for Clk_period;
		Addr <=  "00010011001010";
		Trees_din <= x"08001704";
		wait for Clk_period;
		Addr <=  "00010011001011";
		Trees_din <= x"004913f9";
		wait for Clk_period;
		Addr <=  "00010011001100";
		Trees_din <= x"000e13f9";
		wait for Clk_period;
		Addr <=  "00010011001101";
		Trees_din <= x"1d005004";
		wait for Clk_period;
		Addr <=  "00010011001110";
		Trees_din <= x"009613f9";
		wait for Clk_period;
		Addr <=  "00010011001111";
		Trees_din <= x"ffa713f9";
		wait for Clk_period;
		Addr <=  "00010011010000";
		Trees_din <= x"1900ac10";
		wait for Clk_period;
		Addr <=  "00010011010001";
		Trees_din <= x"010ea208";
		wait for Clk_period;
		Addr <=  "00010011010010";
		Trees_din <= x"06f86a04";
		wait for Clk_period;
		Addr <=  "00010011010011";
		Trees_din <= x"00a913f9";
		wait for Clk_period;
		Addr <=  "00010011010100";
		Trees_din <= x"000f13f9";
		wait for Clk_period;
		Addr <=  "00010011010101";
		Trees_din <= x"0f00a304";
		wait for Clk_period;
		Addr <=  "00010011010110";
		Trees_din <= x"ff8613f9";
		wait for Clk_period;
		Addr <=  "00010011010111";
		Trees_din <= x"005213f9";
		wait for Clk_period;
		Addr <=  "00010011011000";
		Trees_din <= x"07005208";
		wait for Clk_period;
		Addr <=  "00010011011001";
		Trees_din <= x"08005e04";
		wait for Clk_period;
		Addr <=  "00010011011010";
		Trees_din <= x"ffcd13f9";
		wait for Clk_period;
		Addr <=  "00010011011011";
		Trees_din <= x"006413f9";
		wait for Clk_period;
		Addr <=  "00010011011100";
		Trees_din <= x"1900b904";
		wait for Clk_period;
		Addr <=  "00010011011101";
		Trees_din <= x"ffc713f9";
		wait for Clk_period;
		Addr <=  "00010011011110";
		Trees_din <= x"00ba13f9";
		wait for Clk_period;
		Addr <=  "00010011011111";
		Trees_din <= x"010d4f20";
		wait for Clk_period;
		Addr <=  "00010011100000";
		Trees_din <= x"0a07cb18";
		wait for Clk_period;
		Addr <=  "00010011100001";
		Trees_din <= x"0d000008";
		wait for Clk_period;
		Addr <=  "00010011100010";
		Trees_din <= x"1c003204";
		wait for Clk_period;
		Addr <=  "00010011100011";
		Trees_din <= x"ffb913f9";
		wait for Clk_period;
		Addr <=  "00010011100100";
		Trees_din <= x"007313f9";
		wait for Clk_period;
		Addr <=  "00010011100101";
		Trees_din <= x"1f000c08";
		wait for Clk_period;
		Addr <=  "00010011100110";
		Trees_din <= x"21000004";
		wait for Clk_period;
		Addr <=  "00010011100111";
		Trees_din <= x"009c13f9";
		wait for Clk_period;
		Addr <=  "00010011101000";
		Trees_din <= x"005a13f9";
		wait for Clk_period;
		Addr <=  "00010011101001";
		Trees_din <= x"01065e04";
		wait for Clk_period;
		Addr <=  "00010011101010";
		Trees_din <= x"007b13f9";
		wait for Clk_period;
		Addr <=  "00010011101011";
		Trees_din <= x"ffb713f9";
		wait for Clk_period;
		Addr <=  "00010011101100";
		Trees_din <= x"05fc5204";
		wait for Clk_period;
		Addr <=  "00010011101101";
		Trees_din <= x"005613f9";
		wait for Clk_period;
		Addr <=  "00010011101110";
		Trees_din <= x"ffc513f9";
		wait for Clk_period;
		Addr <=  "00010011101111";
		Trees_din <= x"1a00c308";
		wait for Clk_period;
		Addr <=  "00010011110000";
		Trees_din <= x"0801d404";
		wait for Clk_period;
		Addr <=  "00010011110001";
		Trees_din <= x"009213f9";
		wait for Clk_period;
		Addr <=  "00010011110010";
		Trees_din <= x"000013f9";
		wait for Clk_period;
		Addr <=  "00010011110011";
		Trees_din <= x"1e00660c";
		wait for Clk_period;
		Addr <=  "00010011110100";
		Trees_din <= x"00192f08";
		wait for Clk_period;
		Addr <=  "00010011110101";
		Trees_din <= x"0d01a304";
		wait for Clk_period;
		Addr <=  "00010011110110";
		Trees_din <= x"ffbc13f9";
		wait for Clk_period;
		Addr <=  "00010011110111";
		Trees_din <= x"007613f9";
		wait for Clk_period;
		Addr <=  "00010011111000";
		Trees_din <= x"008c13f9";
		wait for Clk_period;
		Addr <=  "00010011111001";
		Trees_din <= x"17000004";
		wait for Clk_period;
		Addr <=  "00010011111010";
		Trees_din <= x"006213f9";
		wait for Clk_period;
		Addr <=  "00010011111011";
		Trees_din <= x"001be904";
		wait for Clk_period;
		Addr <=  "00010011111100";
		Trees_din <= x"ff2d13f9";
		wait for Clk_period;
		Addr <=  "00010011111101";
		Trees_din <= x"fff613f9";
		wait for Clk_period;
		Addr <=  "00010011111110";
		Trees_din <= x"00167668";
		wait for Clk_period;
		Addr <=  "00010011111111";
		Trees_din <= x"0004c628";
		wait for Clk_period;
		Addr <=  "00010100000000";
		Trees_din <= x"0205f220";
		wait for Clk_period;
		Addr <=  "00010100000001";
		Trees_din <= x"02037010";
		wait for Clk_period;
		Addr <=  "00010100000010";
		Trees_din <= x"0f036808";
		wait for Clk_period;
		Addr <=  "00010100000011";
		Trees_din <= x"1a010504";
		wait for Clk_period;
		Addr <=  "00010100000100";
		Trees_din <= x"ffad1535";
		wait for Clk_period;
		Addr <=  "00010100000101";
		Trees_din <= x"00551535";
		wait for Clk_period;
		Addr <=  "00010100000110";
		Trees_din <= x"07005804";
		wait for Clk_period;
		Addr <=  "00010100000111";
		Trees_din <= x"00931535";
		wait for Clk_period;
		Addr <=  "00010100001000";
		Trees_din <= x"ff891535";
		wait for Clk_period;
		Addr <=  "00010100001001";
		Trees_din <= x"0f007f08";
		wait for Clk_period;
		Addr <=  "00010100001010";
		Trees_din <= x"04025d04";
		wait for Clk_period;
		Addr <=  "00010100001011";
		Trees_din <= x"001f1535";
		wait for Clk_period;
		Addr <=  "00010100001100";
		Trees_din <= x"00fc1535";
		wait for Clk_period;
		Addr <=  "00010100001101";
		Trees_din <= x"1102eb04";
		wait for Clk_period;
		Addr <=  "00010100001110";
		Trees_din <= x"ff7e1535";
		wait for Clk_period;
		Addr <=  "00010100001111";
		Trees_din <= x"00a41535";
		wait for Clk_period;
		Addr <=  "00010100010000";
		Trees_din <= x"0bf94004";
		wait for Clk_period;
		Addr <=  "00010100010001";
		Trees_din <= x"00271535";
		wait for Clk_period;
		Addr <=  "00010100010010";
		Trees_din <= x"ff691535";
		wait for Clk_period;
		Addr <=  "00010100010011";
		Trees_din <= x"06f37f20";
		wait for Clk_period;
		Addr <=  "00010100010100";
		Trees_din <= x"0203d010";
		wait for Clk_period;
		Addr <=  "00010100010101";
		Trees_din <= x"0f03bf08";
		wait for Clk_period;
		Addr <=  "00010100010110";
		Trees_din <= x"0a03a304";
		wait for Clk_period;
		Addr <=  "00010100010111";
		Trees_din <= x"00b41535";
		wait for Clk_period;
		Addr <=  "00010100011000";
		Trees_din <= x"ffd51535";
		wait for Clk_period;
		Addr <=  "00010100011001";
		Trees_din <= x"05fa1004";
		wait for Clk_period;
		Addr <=  "00010100011010";
		Trees_din <= x"00691535";
		wait for Clk_period;
		Addr <=  "00010100011011";
		Trees_din <= x"ff901535";
		wait for Clk_period;
		Addr <=  "00010100011100";
		Trees_din <= x"0e012008";
		wait for Clk_period;
		Addr <=  "00010100011101";
		Trees_din <= x"1c004204";
		wait for Clk_period;
		Addr <=  "00010100011110";
		Trees_din <= x"007b1535";
		wait for Clk_period;
		Addr <=  "00010100011111";
		Trees_din <= x"ffc31535";
		wait for Clk_period;
		Addr <=  "00010100100000";
		Trees_din <= x"03fee204";
		wait for Clk_period;
		Addr <=  "00010100100001";
		Trees_din <= x"ffc91535";
		wait for Clk_period;
		Addr <=  "00010100100010";
		Trees_din <= x"00b51535";
		wait for Clk_period;
		Addr <=  "00010100100011";
		Trees_din <= x"0c036410";
		wait for Clk_period;
		Addr <=  "00010100100100";
		Trees_din <= x"1f000008";
		wait for Clk_period;
		Addr <=  "00010100100101";
		Trees_din <= x"06f45804";
		wait for Clk_period;
		Addr <=  "00010100100110";
		Trees_din <= x"ffc51535";
		wait for Clk_period;
		Addr <=  "00010100100111";
		Trees_din <= x"00191535";
		wait for Clk_period;
		Addr <=  "00010100101000";
		Trees_din <= x"0b028804";
		wait for Clk_period;
		Addr <=  "00010100101001";
		Trees_din <= x"00861535";
		wait for Clk_period;
		Addr <=  "00010100101010";
		Trees_din <= x"00131535";
		wait for Clk_period;
		Addr <=  "00010100101011";
		Trees_din <= x"0d004d08";
		wait for Clk_period;
		Addr <=  "00010100101100";
		Trees_din <= x"1d004a04";
		wait for Clk_period;
		Addr <=  "00010100101101";
		Trees_din <= x"009d1535";
		wait for Clk_period;
		Addr <=  "00010100101110";
		Trees_din <= x"001f1535";
		wait for Clk_period;
		Addr <=  "00010100101111";
		Trees_din <= x"05fcf804";
		wait for Clk_period;
		Addr <=  "00010100110000";
		Trees_din <= x"ffb51535";
		wait for Clk_period;
		Addr <=  "00010100110001";
		Trees_din <= x"00221535";
		wait for Clk_period;
		Addr <=  "00010100110010";
		Trees_din <= x"010d4f18";
		wait for Clk_period;
		Addr <=  "00010100110011";
		Trees_din <= x"0f03d40c";
		wait for Clk_period;
		Addr <=  "00010100110100";
		Trees_din <= x"21000004";
		wait for Clk_period;
		Addr <=  "00010100110101";
		Trees_din <= x"009b1535";
		wait for Clk_period;
		Addr <=  "00010100110110";
		Trees_din <= x"19008e04";
		wait for Clk_period;
		Addr <=  "00010100110111";
		Trees_din <= x"ffbe1535";
		wait for Clk_period;
		Addr <=  "00010100111000";
		Trees_din <= x"00781535";
		wait for Clk_period;
		Addr <=  "00010100111001";
		Trees_din <= x"1c003108";
		wait for Clk_period;
		Addr <=  "00010100111010";
		Trees_din <= x"10027a04";
		wait for Clk_period;
		Addr <=  "00010100111011";
		Trees_din <= x"ff041535";
		wait for Clk_period;
		Addr <=  "00010100111100";
		Trees_din <= x"005a1535";
		wait for Clk_period;
		Addr <=  "00010100111101";
		Trees_din <= x"00901535";
		wait for Clk_period;
		Addr <=  "00010100111110";
		Trees_din <= x"1a00c308";
		wait for Clk_period;
		Addr <=  "00010100111111";
		Trees_din <= x"0801d404";
		wait for Clk_period;
		Addr <=  "00010101000000";
		Trees_din <= x"008e1535";
		wait for Clk_period;
		Addr <=  "00010101000001";
		Trees_din <= x"fffe1535";
		wait for Clk_period;
		Addr <=  "00010101000010";
		Trees_din <= x"1e00660c";
		wait for Clk_period;
		Addr <=  "00010101000011";
		Trees_din <= x"00192f08";
		wait for Clk_period;
		Addr <=  "00010101000100";
		Trees_din <= x"0d01a304";
		wait for Clk_period;
		Addr <=  "00010101000101";
		Trees_din <= x"ffc41535";
		wait for Clk_period;
		Addr <=  "00010101000110";
		Trees_din <= x"00701535";
		wait for Clk_period;
		Addr <=  "00010101000111";
		Trees_din <= x"00871535";
		wait for Clk_period;
		Addr <=  "00010101001000";
		Trees_din <= x"17000004";
		wait for Clk_period;
		Addr <=  "00010101001001";
		Trees_din <= x"005c1535";
		wait for Clk_period;
		Addr <=  "00010101001010";
		Trees_din <= x"13fdc604";
		wait for Clk_period;
		Addr <=  "00010101001011";
		Trees_din <= x"001c1535";
		wait for Clk_period;
		Addr <=  "00010101001100";
		Trees_din <= x"ff551535";
		wait for Clk_period;
		Addr <=  "00010101001101";
		Trees_din <= x"00167670";
		wait for Clk_period;
		Addr <=  "00010101001110";
		Trees_din <= x"00079038";
		wait for Clk_period;
		Addr <=  "00010101001111";
		Trees_din <= x"13ffd51c";
		wait for Clk_period;
		Addr <=  "00010101010000";
		Trees_din <= x"0103410c";
		wait for Clk_period;
		Addr <=  "00010101010001";
		Trees_din <= x"11fed304";
		wait for Clk_period;
		Addr <=  "00010101010010";
		Trees_din <= x"ff711689";
		wait for Clk_period;
		Addr <=  "00010101010011";
		Trees_din <= x"00019004";
		wait for Clk_period;
		Addr <=  "00010101010100";
		Trees_din <= x"ffbd1689";
		wait for Clk_period;
		Addr <=  "00010101010101";
		Trees_din <= x"00371689";
		wait for Clk_period;
		Addr <=  "00010101010110";
		Trees_din <= x"04065f08";
		wait for Clk_period;
		Addr <=  "00010101010111";
		Trees_din <= x"07005d04";
		wait for Clk_period;
		Addr <=  "00010101011000";
		Trees_din <= x"ff7c1689";
		wait for Clk_period;
		Addr <=  "00010101011001";
		Trees_din <= x"004a1689";
		wait for Clk_period;
		Addr <=  "00010101011010";
		Trees_din <= x"0b04af04";
		wait for Clk_period;
		Addr <=  "00010101011011";
		Trees_din <= x"ffc31689";
		wait for Clk_period;
		Addr <=  "00010101011100";
		Trees_din <= x"00d21689";
		wait for Clk_period;
		Addr <=  "00010101011101";
		Trees_din <= x"07005610";
		wait for Clk_period;
		Addr <=  "00010101011110";
		Trees_din <= x"0bfa3808";
		wait for Clk_period;
		Addr <=  "00010101011111";
		Trees_din <= x"05fdf604";
		wait for Clk_period;
		Addr <=  "00010101100000";
		Trees_din <= x"00dc1689";
		wait for Clk_period;
		Addr <=  "00010101100001";
		Trees_din <= x"00051689";
		wait for Clk_period;
		Addr <=  "00010101100010";
		Trees_din <= x"0d012d04";
		wait for Clk_period;
		Addr <=  "00010101100011";
		Trees_din <= x"007c1689";
		wait for Clk_period;
		Addr <=  "00010101100100";
		Trees_din <= x"ffbe1689";
		wait for Clk_period;
		Addr <=  "00010101100101";
		Trees_din <= x"05fd1d04";
		wait for Clk_period;
		Addr <=  "00010101100110";
		Trees_din <= x"ff6b1689";
		wait for Clk_period;
		Addr <=  "00010101100111";
		Trees_din <= x"0800e704";
		wait for Clk_period;
		Addr <=  "00010101101000";
		Trees_din <= x"008d1689";
		wait for Clk_period;
		Addr <=  "00010101101001";
		Trees_din <= x"ff8f1689";
		wait for Clk_period;
		Addr <=  "00010101101010";
		Trees_din <= x"04ff5720";
		wait for Clk_period;
		Addr <=  "00010101101011";
		Trees_din <= x"07005b10";
		wait for Clk_period;
		Addr <=  "00010101101100";
		Trees_din <= x"0bf8e908";
		wait for Clk_period;
		Addr <=  "00010101101101";
		Trees_din <= x"1b003304";
		wait for Clk_period;
		Addr <=  "00010101101110";
		Trees_din <= x"00071689";
		wait for Clk_period;
		Addr <=  "00010101101111";
		Trees_din <= x"00af1689";
		wait for Clk_period;
		Addr <=  "00010101110000";
		Trees_din <= x"0c033104";
		wait for Clk_period;
		Addr <=  "00010101110001";
		Trees_din <= x"001c1689";
		wait for Clk_period;
		Addr <=  "00010101110010";
		Trees_din <= x"ffe11689";
		wait for Clk_period;
		Addr <=  "00010101110011";
		Trees_din <= x"0105f908";
		wait for Clk_period;
		Addr <=  "00010101110100";
		Trees_din <= x"01fd2104";
		wait for Clk_period;
		Addr <=  "00010101110101";
		Trees_din <= x"ff9e1689";
		wait for Clk_period;
		Addr <=  "00010101110110";
		Trees_din <= x"00541689";
		wait for Clk_period;
		Addr <=  "00010101110111";
		Trees_din <= x"0f010304";
		wait for Clk_period;
		Addr <=  "00010101111000";
		Trees_din <= x"ffff1689";
		wait for Clk_period;
		Addr <=  "00010101111001";
		Trees_din <= x"ff7d1689";
		wait for Clk_period;
		Addr <=  "00010101111010";
		Trees_din <= x"1c004d10";
		wait for Clk_period;
		Addr <=  "00010101111011";
		Trees_din <= x"08000b08";
		wait for Clk_period;
		Addr <=  "00010101111100";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00010101111101";
		Trees_din <= x"ff341689";
		wait for Clk_period;
		Addr <=  "00010101111110";
		Trees_din <= x"00321689";
		wait for Clk_period;
		Addr <=  "00010101111111";
		Trees_din <= x"05fe3104";
		wait for Clk_period;
		Addr <=  "00010110000000";
		Trees_din <= x"00761689";
		wait for Clk_period;
		Addr <=  "00010110000001";
		Trees_din <= x"ffc71689";
		wait for Clk_period;
		Addr <=  "00010110000010";
		Trees_din <= x"0c013004";
		wait for Clk_period;
		Addr <=  "00010110000011";
		Trees_din <= x"fffe1689";
		wait for Clk_period;
		Addr <=  "00010110000100";
		Trees_din <= x"ff531689";
		wait for Clk_period;
		Addr <=  "00010110000101";
		Trees_din <= x"010d4f18";
		wait for Clk_period;
		Addr <=  "00010110000110";
		Trees_din <= x"0f03d40c";
		wait for Clk_period;
		Addr <=  "00010110000111";
		Trees_din <= x"21000004";
		wait for Clk_period;
		Addr <=  "00010110001000";
		Trees_din <= x"009a1689";
		wait for Clk_period;
		Addr <=  "00010110001001";
		Trees_din <= x"11028104";
		wait for Clk_period;
		Addr <=  "00010110001010";
		Trees_din <= x"00711689";
		wait for Clk_period;
		Addr <=  "00010110001011";
		Trees_din <= x"ffb61689";
		wait for Clk_period;
		Addr <=  "00010110001100";
		Trees_din <= x"1a00dd04";
		wait for Clk_period;
		Addr <=  "00010110001101";
		Trees_din <= x"008d1689";
		wait for Clk_period;
		Addr <=  "00010110001110";
		Trees_din <= x"0102c704";
		wait for Clk_period;
		Addr <=  "00010110001111";
		Trees_din <= x"00541689";
		wait for Clk_period;
		Addr <=  "00010110010000";
		Trees_din <= x"ff191689";
		wait for Clk_period;
		Addr <=  "00010110010001";
		Trees_din <= x"1a00c308";
		wait for Clk_period;
		Addr <=  "00010110010010";
		Trees_din <= x"0801d404";
		wait for Clk_period;
		Addr <=  "00010110010011";
		Trees_din <= x"00891689";
		wait for Clk_period;
		Addr <=  "00010110010100";
		Trees_din <= x"fffe1689";
		wait for Clk_period;
		Addr <=  "00010110010101";
		Trees_din <= x"1e006610";
		wait for Clk_period;
		Addr <=  "00010110010110";
		Trees_din <= x"09005408";
		wait for Clk_period;
		Addr <=  "00010110010111";
		Trees_din <= x"05f75a04";
		wait for Clk_period;
		Addr <=  "00010110011000";
		Trees_din <= x"00101689";
		wait for Clk_period;
		Addr <=  "00010110011001";
		Trees_din <= x"00851689";
		wait for Clk_period;
		Addr <=  "00010110011010";
		Trees_din <= x"1a00db04";
		wait for Clk_period;
		Addr <=  "00010110011011";
		Trees_din <= x"00661689";
		wait for Clk_period;
		Addr <=  "00010110011100";
		Trees_din <= x"ff8f1689";
		wait for Clk_period;
		Addr <=  "00010110011101";
		Trees_din <= x"17000004";
		wait for Clk_period;
		Addr <=  "00010110011110";
		Trees_din <= x"00551689";
		wait for Clk_period;
		Addr <=  "00010110011111";
		Trees_din <= x"001be904";
		wait for Clk_period;
		Addr <=  "00010110100000";
		Trees_din <= x"ff591689";
		wait for Clk_period;
		Addr <=  "00010110100001";
		Trees_din <= x"fffd1689";
		wait for Clk_period;
		Addr <=  "00010110100010";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00010110100011";
		Trees_din <= x"00192f7c";
		wait for Clk_period;
		Addr <=  "00010110100100";
		Trees_din <= x"000b1e3c";
		wait for Clk_period;
		Addr <=  "00010110100101";
		Trees_din <= x"18003d1c";
		wait for Clk_period;
		Addr <=  "00010110100110";
		Trees_din <= x"1c002e10";
		wait for Clk_period;
		Addr <=  "00010110100111";
		Trees_din <= x"08017508";
		wait for Clk_period;
		Addr <=  "00010110101000";
		Trees_din <= x"01018104";
		wait for Clk_period;
		Addr <=  "00010110101001";
		Trees_din <= x"001117c9";
		wait for Clk_period;
		Addr <=  "00010110101010";
		Trees_din <= x"ff8617c9";
		wait for Clk_period;
		Addr <=  "00010110101011";
		Trees_din <= x"0d011504";
		wait for Clk_period;
		Addr <=  "00010110101100";
		Trees_din <= x"ffa817c9";
		wait for Clk_period;
		Addr <=  "00010110101101";
		Trees_din <= x"005117c9";
		wait for Clk_period;
		Addr <=  "00010110101110";
		Trees_din <= x"08001e04";
		wait for Clk_period;
		Addr <=  "00010110101111";
		Trees_din <= x"003b17c9";
		wait for Clk_period;
		Addr <=  "00010110110000";
		Trees_din <= x"07005804";
		wait for Clk_period;
		Addr <=  "00010110110001";
		Trees_din <= x"ff5417c9";
		wait for Clk_period;
		Addr <=  "00010110110010";
		Trees_din <= x"ffd417c9";
		wait for Clk_period;
		Addr <=  "00010110110011";
		Trees_din <= x"19008a10";
		wait for Clk_period;
		Addr <=  "00010110110100";
		Trees_din <= x"04ff7608";
		wait for Clk_period;
		Addr <=  "00010110110101";
		Trees_din <= x"000aa504";
		wait for Clk_period;
		Addr <=  "00010110110110";
		Trees_din <= x"ff6617c9";
		wait for Clk_period;
		Addr <=  "00010110110111";
		Trees_din <= x"002917c9";
		wait for Clk_period;
		Addr <=  "00010110111000";
		Trees_din <= x"05ff8104";
		wait for Clk_period;
		Addr <=  "00010110111001";
		Trees_din <= x"fff017c9";
		wait for Clk_period;
		Addr <=  "00010110111010";
		Trees_din <= x"00bc17c9";
		wait for Clk_period;
		Addr <=  "00010110111011";
		Trees_din <= x"13ff5808";
		wait for Clk_period;
		Addr <=  "00010110111100";
		Trees_din <= x"03fee204";
		wait for Clk_period;
		Addr <=  "00010110111101";
		Trees_din <= x"008617c9";
		wait for Clk_period;
		Addr <=  "00010110111110";
		Trees_din <= x"000017c9";
		wait for Clk_period;
		Addr <=  "00010110111111";
		Trees_din <= x"12021004";
		wait for Clk_period;
		Addr <=  "00010111000000";
		Trees_din <= x"ff8b17c9";
		wait for Clk_period;
		Addr <=  "00010111000001";
		Trees_din <= x"001e17c9";
		wait for Clk_period;
		Addr <=  "00010111000010";
		Trees_din <= x"01082a20";
		wait for Clk_period;
		Addr <=  "00010111000011";
		Trees_din <= x"06f93810";
		wait for Clk_period;
		Addr <=  "00010111000100";
		Trees_din <= x"02045408";
		wait for Clk_period;
		Addr <=  "00010111000101";
		Trees_din <= x"0e052804";
		wait for Clk_period;
		Addr <=  "00010111000110";
		Trees_din <= x"009217c9";
		wait for Clk_period;
		Addr <=  "00010111000111";
		Trees_din <= x"ffe017c9";
		wait for Clk_period;
		Addr <=  "00010111001000";
		Trees_din <= x"0b028804";
		wait for Clk_period;
		Addr <=  "00010111001001";
		Trees_din <= x"004b17c9";
		wait for Clk_period;
		Addr <=  "00010111001010";
		Trees_din <= x"fff117c9";
		wait for Clk_period;
		Addr <=  "00010111001011";
		Trees_din <= x"1400cf08";
		wait for Clk_period;
		Addr <=  "00010111001100";
		Trees_din <= x"11fee804";
		wait for Clk_period;
		Addr <=  "00010111001101";
		Trees_din <= x"002417c9";
		wait for Clk_period;
		Addr <=  "00010111001110";
		Trees_din <= x"009217c9";
		wait for Clk_period;
		Addr <=  "00010111001111";
		Trees_din <= x"1400e004";
		wait for Clk_period;
		Addr <=  "00010111010000";
		Trees_din <= x"fe8317c9";
		wait for Clk_period;
		Addr <=  "00010111010001";
		Trees_din <= x"fff517c9";
		wait for Clk_period;
		Addr <=  "00010111010010";
		Trees_din <= x"08001910";
		wait for Clk_period;
		Addr <=  "00010111010011";
		Trees_din <= x"0b03e308";
		wait for Clk_period;
		Addr <=  "00010111010100";
		Trees_din <= x"0c001f04";
		wait for Clk_period;
		Addr <=  "00010111010101";
		Trees_din <= x"ffa117c9";
		wait for Clk_period;
		Addr <=  "00010111010110";
		Trees_din <= x"00a517c9";
		wait for Clk_period;
		Addr <=  "00010111010111";
		Trees_din <= x"1200c804";
		wait for Clk_period;
		Addr <=  "00010111011000";
		Trees_din <= x"006617c9";
		wait for Clk_period;
		Addr <=  "00010111011001";
		Trees_din <= x"ff9417c9";
		wait for Clk_period;
		Addr <=  "00010111011010";
		Trees_din <= x"05fa5808";
		wait for Clk_period;
		Addr <=  "00010111011011";
		Trees_din <= x"08030104";
		wait for Clk_period;
		Addr <=  "00010111011100";
		Trees_din <= x"002617c9";
		wait for Clk_period;
		Addr <=  "00010111011101";
		Trees_din <= x"ffb017c9";
		wait for Clk_period;
		Addr <=  "00010111011110";
		Trees_din <= x"08007d04";
		wait for Clk_period;
		Addr <=  "00010111011111";
		Trees_din <= x"ff9f17c9";
		wait for Clk_period;
		Addr <=  "00010111100000";
		Trees_din <= x"000517c9";
		wait for Clk_period;
		Addr <=  "00010111100001";
		Trees_din <= x"010ed018";
		wait for Clk_period;
		Addr <=  "00010111100010";
		Trees_din <= x"0d000004";
		wait for Clk_period;
		Addr <=  "00010111100011";
		Trees_din <= x"fff817c9";
		wait for Clk_period;
		Addr <=  "00010111100100";
		Trees_din <= x"1f000c0c";
		wait for Clk_period;
		Addr <=  "00010111100101";
		Trees_din <= x"21000004";
		wait for Clk_period;
		Addr <=  "00010111100110";
		Trees_din <= x"009917c9";
		wait for Clk_period;
		Addr <=  "00010111100111";
		Trees_din <= x"19009204";
		wait for Clk_period;
		Addr <=  "00010111101000";
		Trees_din <= x"ffb717c9";
		wait for Clk_period;
		Addr <=  "00010111101001";
		Trees_din <= x"006617c9";
		wait for Clk_period;
		Addr <=  "00010111101010";
		Trees_din <= x"11025d04";
		wait for Clk_period;
		Addr <=  "00010111101011";
		Trees_din <= x"005e17c9";
		wait for Clk_period;
		Addr <=  "00010111101100";
		Trees_din <= x"ffb917c9";
		wait for Clk_period;
		Addr <=  "00010111101101";
		Trees_din <= x"010fa404";
		wait for Clk_period;
		Addr <=  "00010111101110";
		Trees_din <= x"ffc217c9";
		wait for Clk_period;
		Addr <=  "00010111101111";
		Trees_din <= x"02062104";
		wait for Clk_period;
		Addr <=  "00010111110000";
		Trees_din <= x"007c17c9";
		wait for Clk_period;
		Addr <=  "00010111110001";
		Trees_din <= x"ffe717c9";
		wait for Clk_period;
		Addr <=  "00010111110010";
		Trees_din <= x"00192f54";
		wait for Clk_period;
		Addr <=  "00010111110011";
		Trees_din <= x"0000af18";
		wait for Clk_period;
		Addr <=  "00010111110100";
		Trees_din <= x"09005414";
		wait for Clk_period;
		Addr <=  "00010111110101";
		Trees_din <= x"1101510c";
		wait for Clk_period;
		Addr <=  "00010111110110";
		Trees_din <= x"11010008";
		wait for Clk_period;
		Addr <=  "00010111110111";
		Trees_din <= x"15009104";
		wait for Clk_period;
		Addr <=  "00010111111000";
		Trees_din <= x"002f18bd";
		wait for Clk_period;
		Addr <=  "00010111111001";
		Trees_din <= x"ff9618bd";
		wait for Clk_period;
		Addr <=  "00010111111010";
		Trees_din <= x"011118bd";
		wait for Clk_period;
		Addr <=  "00010111111011";
		Trees_din <= x"02fba504";
		wait for Clk_period;
		Addr <=  "00010111111100";
		Trees_din <= x"004018bd";
		wait for Clk_period;
		Addr <=  "00010111111101";
		Trees_din <= x"ff7e18bd";
		wait for Clk_period;
		Addr <=  "00010111111110";
		Trees_din <= x"ff7318bd";
		wait for Clk_period;
		Addr <=  "00010111111111";
		Trees_din <= x"06f37f20";
		wait for Clk_period;
		Addr <=  "00011000000000";
		Trees_din <= x"0afcf310";
		wait for Clk_period;
		Addr <=  "00011000000001";
		Trees_din <= x"010cd708";
		wait for Clk_period;
		Addr <=  "00011000000010";
		Trees_din <= x"13018c04";
		wait for Clk_period;
		Addr <=  "00011000000011";
		Trees_din <= x"005d18bd";
		wait for Clk_period;
		Addr <=  "00011000000100";
		Trees_din <= x"ff9818bd";
		wait for Clk_period;
		Addr <=  "00011000000101";
		Trees_din <= x"0203d004";
		wait for Clk_period;
		Addr <=  "00011000000110";
		Trees_din <= x"003618bd";
		wait for Clk_period;
		Addr <=  "00011000000111";
		Trees_din <= x"ff7f18bd";
		wait for Clk_period;
		Addr <=  "00011000001000";
		Trees_din <= x"0005c708";
		wait for Clk_period;
		Addr <=  "00011000001001";
		Trees_din <= x"0f000604";
		wait for Clk_period;
		Addr <=  "00011000001010";
		Trees_din <= x"005e18bd";
		wait for Clk_period;
		Addr <=  "00011000001011";
		Trees_din <= x"ff8218bd";
		wait for Clk_period;
		Addr <=  "00011000001100";
		Trees_din <= x"1a00b604";
		wait for Clk_period;
		Addr <=  "00011000001101";
		Trees_din <= x"001818bd";
		wait for Clk_period;
		Addr <=  "00011000001110";
		Trees_din <= x"007b18bd";
		wait for Clk_period;
		Addr <=  "00011000001111";
		Trees_din <= x"0c036410";
		wait for Clk_period;
		Addr <=  "00011000010000";
		Trees_din <= x"00148708";
		wait for Clk_period;
		Addr <=  "00011000010001";
		Trees_din <= x"09005104";
		wait for Clk_period;
		Addr <=  "00011000010010";
		Trees_din <= x"ffe518bd";
		wait for Clk_period;
		Addr <=  "00011000010011";
		Trees_din <= x"001318bd";
		wait for Clk_period;
		Addr <=  "00011000010100";
		Trees_din <= x"03f28904";
		wait for Clk_period;
		Addr <=  "00011000010101";
		Trees_din <= x"ffaa18bd";
		wait for Clk_period;
		Addr <=  "00011000010110";
		Trees_din <= x"005518bd";
		wait for Clk_period;
		Addr <=  "00011000010111";
		Trees_din <= x"1104b708";
		wait for Clk_period;
		Addr <=  "00011000011000";
		Trees_din <= x"1b003204";
		wait for Clk_period;
		Addr <=  "00011000011001";
		Trees_din <= x"003e18bd";
		wait for Clk_period;
		Addr <=  "00011000011010";
		Trees_din <= x"ffc518bd";
		wait for Clk_period;
		Addr <=  "00011000011011";
		Trees_din <= x"008718bd";
		wait for Clk_period;
		Addr <=  "00011000011100";
		Trees_din <= x"010ed018";
		wait for Clk_period;
		Addr <=  "00011000011101";
		Trees_din <= x"0d000004";
		wait for Clk_period;
		Addr <=  "00011000011110";
		Trees_din <= x"fff118bd";
		wait for Clk_period;
		Addr <=  "00011000011111";
		Trees_din <= x"1f000c0c";
		wait for Clk_period;
		Addr <=  "00011000100000";
		Trees_din <= x"21000004";
		wait for Clk_period;
		Addr <=  "00011000100001";
		Trees_din <= x"009818bd";
		wait for Clk_period;
		Addr <=  "00011000100010";
		Trees_din <= x"1b003904";
		wait for Clk_period;
		Addr <=  "00011000100011";
		Trees_din <= x"005e18bd";
		wait for Clk_period;
		Addr <=  "00011000100100";
		Trees_din <= x"ffb518bd";
		wait for Clk_period;
		Addr <=  "00011000100101";
		Trees_din <= x"07005604";
		wait for Clk_period;
		Addr <=  "00011000100110";
		Trees_din <= x"005718bd";
		wait for Clk_period;
		Addr <=  "00011000100111";
		Trees_din <= x"ffba18bd";
		wait for Clk_period;
		Addr <=  "00011000101000";
		Trees_din <= x"1d004304";
		wait for Clk_period;
		Addr <=  "00011000101001";
		Trees_din <= x"007518bd";
		wait for Clk_period;
		Addr <=  "00011000101010";
		Trees_din <= x"15009608";
		wait for Clk_period;
		Addr <=  "00011000101011";
		Trees_din <= x"02016004";
		wait for Clk_period;
		Addr <=  "00011000101100";
		Trees_din <= x"ffc718bd";
		wait for Clk_period;
		Addr <=  "00011000101101";
		Trees_din <= x"005d18bd";
		wait for Clk_period;
		Addr <=  "00011000101110";
		Trees_din <= x"ff8f18bd";
		wait for Clk_period;
		Addr <=  "00011000101111";
		Trees_din <= x"00192f68";
		wait for Clk_period;
		Addr <=  "00011000110000";
		Trees_din <= x"0003aa30";
		wait for Clk_period;
		Addr <=  "00011000110001";
		Trees_din <= x"0900541c";
		wait for Clk_period;
		Addr <=  "00011000110010";
		Trees_din <= x"0900500c";
		wait for Clk_period;
		Addr <=  "00011000110011";
		Trees_din <= x"0d001004";
		wait for Clk_period;
		Addr <=  "00011000110100";
		Trees_din <= x"005819c9";
		wait for Clk_period;
		Addr <=  "00011000110101";
		Trees_din <= x"10f99904";
		wait for Clk_period;
		Addr <=  "00011000110110";
		Trees_din <= x"ffee19c9";
		wait for Clk_period;
		Addr <=  "00011000110111";
		Trees_din <= x"ff7619c9";
		wait for Clk_period;
		Addr <=  "00011000111000";
		Trees_din <= x"1e006108";
		wait for Clk_period;
		Addr <=  "00011000111001";
		Trees_din <= x"18003104";
		wait for Clk_period;
		Addr <=  "00011000111010";
		Trees_din <= x"005d19c9";
		wait for Clk_period;
		Addr <=  "00011000111011";
		Trees_din <= x"ff8d19c9";
		wait for Clk_period;
		Addr <=  "00011000111100";
		Trees_din <= x"10041004";
		wait for Clk_period;
		Addr <=  "00011000111101";
		Trees_din <= x"00c919c9";
		wait for Clk_period;
		Addr <=  "00011000111110";
		Trees_din <= x"ff9f19c9";
		wait for Clk_period;
		Addr <=  "00011000111111";
		Trees_din <= x"0bf94008";
		wait for Clk_period;
		Addr <=  "00011001000000";
		Trees_din <= x"1b004304";
		wait for Clk_period;
		Addr <=  "00011001000001";
		Trees_din <= x"ffef19c9";
		wait for Clk_period;
		Addr <=  "00011001000010";
		Trees_din <= x"00a619c9";
		wait for Clk_period;
		Addr <=  "00011001000011";
		Trees_din <= x"01fd7808";
		wait for Clk_period;
		Addr <=  "00011001000100";
		Trees_din <= x"00019004";
		wait for Clk_period;
		Addr <=  "00011001000101";
		Trees_din <= x"ff8919c9";
		wait for Clk_period;
		Addr <=  "00011001000110";
		Trees_din <= x"003319c9";
		wait for Clk_period;
		Addr <=  "00011001000111";
		Trees_din <= x"ff6b19c9";
		wait for Clk_period;
		Addr <=  "00011001001000";
		Trees_din <= x"02fdcd18";
		wait for Clk_period;
		Addr <=  "00011001001001";
		Trees_din <= x"00054508";
		wait for Clk_period;
		Addr <=  "00011001001010";
		Trees_din <= x"12008804";
		wait for Clk_period;
		Addr <=  "00011001001011";
		Trees_din <= x"007a19c9";
		wait for Clk_period;
		Addr <=  "00011001001100";
		Trees_din <= x"ff8319c9";
		wait for Clk_period;
		Addr <=  "00011001001101";
		Trees_din <= x"0f02d608";
		wait for Clk_period;
		Addr <=  "00011001001110";
		Trees_din <= x"02fc0c04";
		wait for Clk_period;
		Addr <=  "00011001001111";
		Trees_din <= x"fff519c9";
		wait for Clk_period;
		Addr <=  "00011001010000";
		Trees_din <= x"00a019c9";
		wait for Clk_period;
		Addr <=  "00011001010001";
		Trees_din <= x"10028504";
		wait for Clk_period;
		Addr <=  "00011001010010";
		Trees_din <= x"ff9d19c9";
		wait for Clk_period;
		Addr <=  "00011001010011";
		Trees_din <= x"003a19c9";
		wait for Clk_period;
		Addr <=  "00011001010100";
		Trees_din <= x"06f37f10";
		wait for Clk_period;
		Addr <=  "00011001010101";
		Trees_din <= x"0005c708";
		wait for Clk_period;
		Addr <=  "00011001010110";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00011001010111";
		Trees_din <= x"001519c9";
		wait for Clk_period;
		Addr <=  "00011001011000";
		Trees_din <= x"ff6f19c9";
		wait for Clk_period;
		Addr <=  "00011001011001";
		Trees_din <= x"03ff5404";
		wait for Clk_period;
		Addr <=  "00011001011010";
		Trees_din <= x"002819c9";
		wait for Clk_period;
		Addr <=  "00011001011011";
		Trees_din <= x"00a619c9";
		wait for Clk_period;
		Addr <=  "00011001011100";
		Trees_din <= x"09005808";
		wait for Clk_period;
		Addr <=  "00011001011101";
		Trees_din <= x"1200fb04";
		wait for Clk_period;
		Addr <=  "00011001011110";
		Trees_din <= x"ffdd19c9";
		wait for Clk_period;
		Addr <=  "00011001011111";
		Trees_din <= x"000919c9";
		wait for Clk_period;
		Addr <=  "00011001100000";
		Trees_din <= x"16018d04";
		wait for Clk_period;
		Addr <=  "00011001100001";
		Trees_din <= x"fff619c9";
		wait for Clk_period;
		Addr <=  "00011001100010";
		Trees_din <= x"004919c9";
		wait for Clk_period;
		Addr <=  "00011001100011";
		Trees_din <= x"01079608";
		wait for Clk_period;
		Addr <=  "00011001100100";
		Trees_din <= x"0d000004";
		wait for Clk_period;
		Addr <=  "00011001100101";
		Trees_din <= x"ffd819c9";
		wait for Clk_period;
		Addr <=  "00011001100110";
		Trees_din <= x"009619c9";
		wait for Clk_period;
		Addr <=  "00011001100111";
		Trees_din <= x"11045114";
		wait for Clk_period;
		Addr <=  "00011001101000";
		Trees_din <= x"0f03d00c";
		wait for Clk_period;
		Addr <=  "00011001101001";
		Trees_din <= x"1703dc08";
		wait for Clk_period;
		Addr <=  "00011001101010";
		Trees_din <= x"0112d604";
		wait for Clk_period;
		Addr <=  "00011001101011";
		Trees_din <= x"008c19c9";
		wait for Clk_period;
		Addr <=  "00011001101100";
		Trees_din <= x"001719c9";
		wait for Clk_period;
		Addr <=  "00011001101101";
		Trees_din <= x"ffe219c9";
		wait for Clk_period;
		Addr <=  "00011001101110";
		Trees_din <= x"16004204";
		wait for Clk_period;
		Addr <=  "00011001101111";
		Trees_din <= x"006019c9";
		wait for Clk_period;
		Addr <=  "00011001110000";
		Trees_din <= x"ff5b19c9";
		wait for Clk_period;
		Addr <=  "00011001110001";
		Trees_din <= x"ffa919c9";
		wait for Clk_period;
		Addr <=  "00011001110010";
		Trees_din <= x"00192f64";
		wait for Clk_period;
		Addr <=  "00011001110011";
		Trees_din <= x"000b1e34";
		wait for Clk_period;
		Addr <=  "00011001110100";
		Trees_din <= x"06f6a514";
		wait for Clk_period;
		Addr <=  "00011001110101";
		Trees_din <= x"020cbe10";
		wait for Clk_period;
		Addr <=  "00011001110110";
		Trees_din <= x"11fed308";
		wait for Clk_period;
		Addr <=  "00011001110111";
		Trees_din <= x"02038004";
		wait for Clk_period;
		Addr <=  "00011001111000";
		Trees_din <= x"00011ac5";
		wait for Clk_period;
		Addr <=  "00011001111001";
		Trees_din <= x"ff661ac5";
		wait for Clk_period;
		Addr <=  "00011001111010";
		Trees_din <= x"0f016e04";
		wait for Clk_period;
		Addr <=  "00011001111011";
		Trees_din <= x"00431ac5";
		wait for Clk_period;
		Addr <=  "00011001111100";
		Trees_din <= x"ffee1ac5";
		wait for Clk_period;
		Addr <=  "00011001111101";
		Trees_din <= x"ff761ac5";
		wait for Clk_period;
		Addr <=  "00011001111110";
		Trees_din <= x"0c017210";
		wait for Clk_period;
		Addr <=  "00011001111111";
		Trees_din <= x"1603fc08";
		wait for Clk_period;
		Addr <=  "00011010000000";
		Trees_din <= x"1a00b104";
		wait for Clk_period;
		Addr <=  "00011010000001";
		Trees_din <= x"ffef1ac5";
		wait for Clk_period;
		Addr <=  "00011010000010";
		Trees_din <= x"ff651ac5";
		wait for Clk_period;
		Addr <=  "00011010000011";
		Trees_din <= x"01024404";
		wait for Clk_period;
		Addr <=  "00011010000100";
		Trees_din <= x"00681ac5";
		wait for Clk_period;
		Addr <=  "00011010000101";
		Trees_din <= x"ffae1ac5";
		wait for Clk_period;
		Addr <=  "00011010000110";
		Trees_din <= x"0f01c208";
		wait for Clk_period;
		Addr <=  "00011010000111";
		Trees_din <= x"13f90804";
		wait for Clk_period;
		Addr <=  "00011010001000";
		Trees_din <= x"00571ac5";
		wait for Clk_period;
		Addr <=  "00011010001001";
		Trees_din <= x"ffb51ac5";
		wait for Clk_period;
		Addr <=  "00011010001010";
		Trees_din <= x"06f76004";
		wait for Clk_period;
		Addr <=  "00011010001011";
		Trees_din <= x"ff9d1ac5";
		wait for Clk_period;
		Addr <=  "00011010001100";
		Trees_din <= x"006d1ac5";
		wait for Clk_period;
		Addr <=  "00011010001101";
		Trees_din <= x"18003610";
		wait for Clk_period;
		Addr <=  "00011010001110";
		Trees_din <= x"020db70c";
		wait for Clk_period;
		Addr <=  "00011010001111";
		Trees_din <= x"1006a808";
		wait for Clk_period;
		Addr <=  "00011010010000";
		Trees_din <= x"14008c04";
		wait for Clk_period;
		Addr <=  "00011010010001";
		Trees_din <= x"fffe1ac5";
		wait for Clk_period;
		Addr <=  "00011010010010";
		Trees_din <= x"00861ac5";
		wait for Clk_period;
		Addr <=  "00011010010011";
		Trees_din <= x"ffac1ac5";
		wait for Clk_period;
		Addr <=  "00011010010100";
		Trees_din <= x"ff841ac5";
		wait for Clk_period;
		Addr <=  "00011010010101";
		Trees_din <= x"1e005b10";
		wait for Clk_period;
		Addr <=  "00011010010110";
		Trees_din <= x"0202e708";
		wait for Clk_period;
		Addr <=  "00011010010111";
		Trees_din <= x"1e005604";
		wait for Clk_period;
		Addr <=  "00011010011000";
		Trees_din <= x"ffa51ac5";
		wait for Clk_period;
		Addr <=  "00011010011001";
		Trees_din <= x"005e1ac5";
		wait for Clk_period;
		Addr <=  "00011010011010";
		Trees_din <= x"05f92804";
		wait for Clk_period;
		Addr <=  "00011010011011";
		Trees_din <= x"001c1ac5";
		wait for Clk_period;
		Addr <=  "00011010011100";
		Trees_din <= x"ff5a1ac5";
		wait for Clk_period;
		Addr <=  "00011010011101";
		Trees_din <= x"0afafe08";
		wait for Clk_period;
		Addr <=  "00011010011110";
		Trees_din <= x"11009004";
		wait for Clk_period;
		Addr <=  "00011010011111";
		Trees_din <= x"007e1ac5";
		wait for Clk_period;
		Addr <=  "00011010100000";
		Trees_din <= x"ffd91ac5";
		wait for Clk_period;
		Addr <=  "00011010100001";
		Trees_din <= x"15008504";
		wait for Clk_period;
		Addr <=  "00011010100010";
		Trees_din <= x"00551ac5";
		wait for Clk_period;
		Addr <=  "00011010100011";
		Trees_din <= x"00141ac5";
		wait for Clk_period;
		Addr <=  "00011010100100";
		Trees_din <= x"01079608";
		wait for Clk_period;
		Addr <=  "00011010100101";
		Trees_din <= x"13f83104";
		wait for Clk_period;
		Addr <=  "00011010100110";
		Trees_din <= x"ffca1ac5";
		wait for Clk_period;
		Addr <=  "00011010100111";
		Trees_din <= x"00941ac5";
		wait for Clk_period;
		Addr <=  "00011010101000";
		Trees_din <= x"13ffb908";
		wait for Clk_period;
		Addr <=  "00011010101001";
		Trees_din <= x"06f26204";
		wait for Clk_period;
		Addr <=  "00011010101010";
		Trees_din <= x"ffeb1ac5";
		wait for Clk_period;
		Addr <=  "00011010101011";
		Trees_din <= x"00871ac5";
		wait for Clk_period;
		Addr <=  "00011010101100";
		Trees_din <= x"0201e308";
		wait for Clk_period;
		Addr <=  "00011010101101";
		Trees_din <= x"0afc9804";
		wait for Clk_period;
		Addr <=  "00011010101110";
		Trees_din <= x"ff011ac5";
		wait for Clk_period;
		Addr <=  "00011010101111";
		Trees_din <= x"00101ac5";
		wait for Clk_period;
		Addr <=  "00011010110000";
		Trees_din <= x"00721ac5";
		wait for Clk_period;
		Addr <=  "00011010110001";
		Trees_din <= x"00192f34";
		wait for Clk_period;
		Addr <=  "00011010110010";
		Trees_din <= x"0000af14";
		wait for Clk_period;
		Addr <=  "00011010110011";
		Trees_din <= x"10f8a608";
		wait for Clk_period;
		Addr <=  "00011010110100";
		Trees_din <= x"12015404";
		wait for Clk_period;
		Addr <=  "00011010110101";
		Trees_din <= x"ffaa1b69";
		wait for Clk_period;
		Addr <=  "00011010110110";
		Trees_din <= x"00c11b69";
		wait for Clk_period;
		Addr <=  "00011010110111";
		Trees_din <= x"08038608";
		wait for Clk_period;
		Addr <=  "00011010111000";
		Trees_din <= x"02fba504";
		wait for Clk_period;
		Addr <=  "00011010111001";
		Trees_din <= x"00171b69";
		wait for Clk_period;
		Addr <=  "00011010111010";
		Trees_din <= x"ff721b69";
		wait for Clk_period;
		Addr <=  "00011010111011";
		Trees_din <= x"004c1b69";
		wait for Clk_period;
		Addr <=  "00011010111100";
		Trees_din <= x"09005e18";
		wait for Clk_period;
		Addr <=  "00011010111101";
		Trees_din <= x"0d03f510";
		wait for Clk_period;
		Addr <=  "00011010111110";
		Trees_din <= x"12fbf708";
		wait for Clk_period;
		Addr <=  "00011010111111";
		Trees_din <= x"04fdef04";
		wait for Clk_period;
		Addr <=  "00011011000000";
		Trees_din <= x"fff41b69";
		wait for Clk_period;
		Addr <=  "00011011000001";
		Trees_din <= x"00ea1b69";
		wait for Clk_period;
		Addr <=  "00011011000010";
		Trees_din <= x"0e06a204";
		wait for Clk_period;
		Addr <=  "00011011000011";
		Trees_din <= x"00031b69";
		wait for Clk_period;
		Addr <=  "00011011000100";
		Trees_din <= x"00831b69";
		wait for Clk_period;
		Addr <=  "00011011000101";
		Trees_din <= x"09005204";
		wait for Clk_period;
		Addr <=  "00011011000110";
		Trees_din <= x"ffd41b69";
		wait for Clk_period;
		Addr <=  "00011011000111";
		Trees_din <= x"00991b69";
		wait for Clk_period;
		Addr <=  "00011011001000";
		Trees_din <= x"01039c04";
		wait for Clk_period;
		Addr <=  "00011011001001";
		Trees_din <= x"ffd01b69";
		wait for Clk_period;
		Addr <=  "00011011001010";
		Trees_din <= x"00a11b69";
		wait for Clk_period;
		Addr <=  "00011011001011";
		Trees_din <= x"06f5b418";
		wait for Clk_period;
		Addr <=  "00011011001100";
		Trees_din <= x"04f5ea08";
		wait for Clk_period;
		Addr <=  "00011011001101";
		Trees_din <= x"0112d604";
		wait for Clk_period;
		Addr <=  "00011011001110";
		Trees_din <= x"00861b69";
		wait for Clk_period;
		Addr <=  "00011011001111";
		Trees_din <= x"00031b69";
		wait for Clk_period;
		Addr <=  "00011011010000";
		Trees_din <= x"0201e308";
		wait for Clk_period;
		Addr <=  "00011011010001";
		Trees_din <= x"06f4df04";
		wait for Clk_period;
		Addr <=  "00011011010010";
		Trees_din <= x"ffee1b69";
		wait for Clk_period;
		Addr <=  "00011011010011";
		Trees_din <= x"fecb1b69";
		wait for Clk_period;
		Addr <=  "00011011010100";
		Trees_din <= x"09004e04";
		wait for Clk_period;
		Addr <=  "00011011010101";
		Trees_din <= x"000d1b69";
		wait for Clk_period;
		Addr <=  "00011011010110";
		Trees_din <= x"00621b69";
		wait for Clk_period;
		Addr <=  "00011011010111";
		Trees_din <= x"1f000c04";
		wait for Clk_period;
		Addr <=  "00011011011000";
		Trees_din <= x"00931b69";
		wait for Clk_period;
		Addr <=  "00011011011001";
		Trees_din <= x"ffdf1b69";
		wait for Clk_period;
		Addr <=  "00011011011010";
		Trees_din <= x"001fa458";
		wait for Clk_period;
		Addr <=  "00011011011011";
		Trees_din <= x"0003aa2c";
		wait for Clk_period;
		Addr <=  "00011011011100";
		Trees_din <= x"07005820";
		wait for Clk_period;
		Addr <=  "00011011011101";
		Trees_din <= x"07005710";
		wait for Clk_period;
		Addr <=  "00011011011110";
		Trees_din <= x"13ffe208";
		wait for Clk_period;
		Addr <=  "00011011011111";
		Trees_din <= x"14003304";
		wait for Clk_period;
		Addr <=  "00011011100000";
		Trees_din <= x"00301c25";
		wait for Clk_period;
		Addr <=  "00011011100001";
		Trees_din <= x"ff801c25";
		wait for Clk_period;
		Addr <=  "00011011100010";
		Trees_din <= x"13fffc04";
		wait for Clk_period;
		Addr <=  "00011011100011";
		Trees_din <= x"00ab1c25";
		wait for Clk_period;
		Addr <=  "00011011100100";
		Trees_din <= x"ffda1c25";
		wait for Clk_period;
		Addr <=  "00011011100101";
		Trees_din <= x"0b028808";
		wait for Clk_period;
		Addr <=  "00011011100110";
		Trees_din <= x"0f004604";
		wait for Clk_period;
		Addr <=  "00011011100111";
		Trees_din <= x"00181c25";
		wait for Clk_period;
		Addr <=  "00011011101000";
		Trees_din <= x"ff921c25";
		wait for Clk_period;
		Addr <=  "00011011101001";
		Trees_din <= x"11013904";
		wait for Clk_period;
		Addr <=  "00011011101010";
		Trees_din <= x"fff31c25";
		wait for Clk_period;
		Addr <=  "00011011101011";
		Trees_din <= x"00fe1c25";
		wait for Clk_period;
		Addr <=  "00011011101100";
		Trees_din <= x"1c002d08";
		wait for Clk_period;
		Addr <=  "00011011101101";
		Trees_din <= x"1500a104";
		wait for Clk_period;
		Addr <=  "00011011101110";
		Trees_din <= x"00591c25";
		wait for Clk_period;
		Addr <=  "00011011101111";
		Trees_din <= x"ffe21c25";
		wait for Clk_period;
		Addr <=  "00011011110000";
		Trees_din <= x"ff731c25";
		wait for Clk_period;
		Addr <=  "00011011110001";
		Trees_din <= x"02fdcd18";
		wait for Clk_period;
		Addr <=  "00011011110010";
		Trees_din <= x"00054508";
		wait for Clk_period;
		Addr <=  "00011011110011";
		Trees_din <= x"12008804";
		wait for Clk_period;
		Addr <=  "00011011110100";
		Trees_din <= x"006b1c25";
		wait for Clk_period;
		Addr <=  "00011011110101";
		Trees_din <= x"ff8e1c25";
		wait for Clk_period;
		Addr <=  "00011011110110";
		Trees_din <= x"0f02d608";
		wait for Clk_period;
		Addr <=  "00011011110111";
		Trees_din <= x"02fc0c04";
		wait for Clk_period;
		Addr <=  "00011011111000";
		Trees_din <= x"fff91c25";
		wait for Clk_period;
		Addr <=  "00011011111001";
		Trees_din <= x"00921c25";
		wait for Clk_period;
		Addr <=  "00011011111010";
		Trees_din <= x"000b9b04";
		wait for Clk_period;
		Addr <=  "00011011111011";
		Trees_din <= x"ffb31c25";
		wait for Clk_period;
		Addr <=  "00011011111100";
		Trees_din <= x"003d1c25";
		wait for Clk_period;
		Addr <=  "00011011111101";
		Trees_din <= x"0306c210";
		wait for Clk_period;
		Addr <=  "00011011111110";
		Trees_din <= x"1900a608";
		wait for Clk_period;
		Addr <=  "00011011111111";
		Trees_din <= x"1b003804";
		wait for Clk_period;
		Addr <=  "00011100000000";
		Trees_din <= x"ffe91c25";
		wait for Clk_period;
		Addr <=  "00011100000001";
		Trees_din <= x"000f1c25";
		wait for Clk_period;
		Addr <=  "00011100000010";
		Trees_din <= x"15009a04";
		wait for Clk_period;
		Addr <=  "00011100000011";
		Trees_din <= x"00851c25";
		wait for Clk_period;
		Addr <=  "00011100000100";
		Trees_din <= x"00111c25";
		wait for Clk_period;
		Addr <=  "00011100000101";
		Trees_din <= x"ff771c25";
		wait for Clk_period;
		Addr <=  "00011100000110";
		Trees_din <= x"1f000c04";
		wait for Clk_period;
		Addr <=  "00011100000111";
		Trees_din <= x"008f1c25";
		wait for Clk_period;
		Addr <=  "00011100001000";
		Trees_din <= x"ffc81c25";
		wait for Clk_period;
		Addr <=  "00011100001001";
		Trees_din <= x"001fa464";
		wait for Clk_period;
		Addr <=  "00011100001010";
		Trees_din <= x"0011923c";
		wait for Clk_period;
		Addr <=  "00011100001011";
		Trees_din <= x"06f79220";
		wait for Clk_period;
		Addr <=  "00011100001100";
		Trees_din <= x"1703e410";
		wait for Clk_period;
		Addr <=  "00011100001101";
		Trees_din <= x"19008308";
		wait for Clk_period;
		Addr <=  "00011100001110";
		Trees_din <= x"1400cc04";
		wait for Clk_period;
		Addr <=  "00011100001111";
		Trees_din <= x"002c1cf9";
		wait for Clk_period;
		Addr <=  "00011100010000";
		Trees_din <= x"ffba1cf9";
		wait for Clk_period;
		Addr <=  "00011100010001";
		Trees_din <= x"1005e404";
		wait for Clk_period;
		Addr <=  "00011100010010";
		Trees_din <= x"00211cf9";
		wait for Clk_period;
		Addr <=  "00011100010011";
		Trees_din <= x"ffac1cf9";
		wait for Clk_period;
		Addr <=  "00011100010100";
		Trees_din <= x"0b03a108";
		wait for Clk_period;
		Addr <=  "00011100010101";
		Trees_din <= x"0afcc504";
		wait for Clk_period;
		Addr <=  "00011100010110";
		Trees_din <= x"ffb21cf9";
		wait for Clk_period;
		Addr <=  "00011100010111";
		Trees_din <= x"00801cf9";
		wait for Clk_period;
		Addr <=  "00011100011000";
		Trees_din <= x"13f85404";
		wait for Clk_period;
		Addr <=  "00011100011001";
		Trees_din <= x"00041cf9";
		wait for Clk_period;
		Addr <=  "00011100011010";
		Trees_din <= x"ff3a1cf9";
		wait for Clk_period;
		Addr <=  "00011100011011";
		Trees_din <= x"0e043e10";
		wait for Clk_period;
		Addr <=  "00011100011100";
		Trees_din <= x"16002008";
		wait for Clk_period;
		Addr <=  "00011100011101";
		Trees_din <= x"1e006e04";
		wait for Clk_period;
		Addr <=  "00011100011110";
		Trees_din <= x"ff381cf9";
		wait for Clk_period;
		Addr <=  "00011100011111";
		Trees_din <= x"00101cf9";
		wait for Clk_period;
		Addr <=  "00011100100000";
		Trees_din <= x"000f9e04";
		wait for Clk_period;
		Addr <=  "00011100100001";
		Trees_din <= x"ffd71cf9";
		wait for Clk_period;
		Addr <=  "00011100100010";
		Trees_din <= x"002f1cf9";
		wait for Clk_period;
		Addr <=  "00011100100011";
		Trees_din <= x"1500a708";
		wait for Clk_period;
		Addr <=  "00011100100100";
		Trees_din <= x"13007e04";
		wait for Clk_period;
		Addr <=  "00011100100101";
		Trees_din <= x"fffb1cf9";
		wait for Clk_period;
		Addr <=  "00011100100110";
		Trees_din <= x"00cf1cf9";
		wait for Clk_period;
		Addr <=  "00011100100111";
		Trees_din <= x"ffaf1cf9";
		wait for Clk_period;
		Addr <=  "00011100101000";
		Trees_din <= x"1500a920";
		wait for Clk_period;
		Addr <=  "00011100101001";
		Trees_din <= x"08015b10";
		wait for Clk_period;
		Addr <=  "00011100101010";
		Trees_din <= x"03f8e608";
		wait for Clk_period;
		Addr <=  "00011100101011";
		Trees_din <= x"03f8a504";
		wait for Clk_period;
		Addr <=  "00011100101100";
		Trees_din <= x"001f1cf9";
		wait for Clk_period;
		Addr <=  "00011100101101";
		Trees_din <= x"ff221cf9";
		wait for Clk_period;
		Addr <=  "00011100101110";
		Trees_din <= x"1b004b04";
		wait for Clk_period;
		Addr <=  "00011100101111";
		Trees_din <= x"00951cf9";
		wait for Clk_period;
		Addr <=  "00011100110000";
		Trees_din <= x"00071cf9";
		wait for Clk_period;
		Addr <=  "00011100110001";
		Trees_din <= x"06f7dd08";
		wait for Clk_period;
		Addr <=  "00011100110010";
		Trees_din <= x"03fa9f04";
		wait for Clk_period;
		Addr <=  "00011100110011";
		Trees_din <= x"ffd81cf9";
		wait for Clk_period;
		Addr <=  "00011100110100";
		Trees_din <= x"feeb1cf9";
		wait for Clk_period;
		Addr <=  "00011100110101";
		Trees_din <= x"0a028704";
		wait for Clk_period;
		Addr <=  "00011100110110";
		Trees_din <= x"00861cf9";
		wait for Clk_period;
		Addr <=  "00011100110111";
		Trees_din <= x"ffcf1cf9";
		wait for Clk_period;
		Addr <=  "00011100111000";
		Trees_din <= x"1d003f04";
		wait for Clk_period;
		Addr <=  "00011100111001";
		Trees_din <= x"00971cf9";
		wait for Clk_period;
		Addr <=  "00011100111010";
		Trees_din <= x"ffb71cf9";
		wait for Clk_period;
		Addr <=  "00011100111011";
		Trees_din <= x"1f000c04";
		wait for Clk_period;
		Addr <=  "00011100111100";
		Trees_din <= x"008d1cf9";
		wait for Clk_period;
		Addr <=  "00011100111101";
		Trees_din <= x"ffd01cf9";
		wait for Clk_period;
		Addr <=  "00011100111110";
		Trees_din <= x"001fa470";
		wait for Clk_period;
		Addr <=  "00011100111111";
		Trees_din <= x"0207143c";
		wait for Clk_period;
		Addr <=  "00011101000000";
		Trees_din <= x"1500921c";
		wait for Clk_period;
		Addr <=  "00011101000001";
		Trees_din <= x"000d9f0c";
		wait for Clk_period;
		Addr <=  "00011101000010";
		Trees_din <= x"10057a08";
		wait for Clk_period;
		Addr <=  "00011101000011";
		Trees_din <= x"1601a604";
		wait for Clk_period;
		Addr <=  "00011101000100";
		Trees_din <= x"ffe01de5";
		wait for Clk_period;
		Addr <=  "00011101000101";
		Trees_din <= x"00361de5";
		wait for Clk_period;
		Addr <=  "00011101000110";
		Trees_din <= x"ff6c1de5";
		wait for Clk_period;
		Addr <=  "00011101000111";
		Trees_din <= x"1c003908";
		wait for Clk_period;
		Addr <=  "00011101001000";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00011101001001";
		Trees_din <= x"ffc51de5";
		wait for Clk_period;
		Addr <=  "00011101001010";
		Trees_din <= x"00b51de5";
		wait for Clk_period;
		Addr <=  "00011101001011";
		Trees_din <= x"1a00ba04";
		wait for Clk_period;
		Addr <=  "00011101001100";
		Trees_din <= x"004a1de5";
		wait for Clk_period;
		Addr <=  "00011101001101";
		Trees_din <= x"ff9c1de5";
		wait for Clk_period;
		Addr <=  "00011101001110";
		Trees_din <= x"1900a310";
		wait for Clk_period;
		Addr <=  "00011101001111";
		Trees_din <= x"06fb8708";
		wait for Clk_period;
		Addr <=  "00011101010000";
		Trees_din <= x"04fb7404";
		wait for Clk_period;
		Addr <=  "00011101010001";
		Trees_din <= x"ffbd1de5";
		wait for Clk_period;
		Addr <=  "00011101010010";
		Trees_din <= x"00011de5";
		wait for Clk_period;
		Addr <=  "00011101010011";
		Trees_din <= x"08001a04";
		wait for Clk_period;
		Addr <=  "00011101010100";
		Trees_din <= x"ff8c1de5";
		wait for Clk_period;
		Addr <=  "00011101010101";
		Trees_din <= x"00671de5";
		wait for Clk_period;
		Addr <=  "00011101010110";
		Trees_din <= x"000fd308";
		wait for Clk_period;
		Addr <=  "00011101010111";
		Trees_din <= x"11fdc204";
		wait for Clk_period;
		Addr <=  "00011101011000";
		Trees_din <= x"ff861de5";
		wait for Clk_period;
		Addr <=  "00011101011001";
		Trees_din <= x"00141de5";
		wait for Clk_period;
		Addr <=  "00011101011010";
		Trees_din <= x"0c01c204";
		wait for Clk_period;
		Addr <=  "00011101011011";
		Trees_din <= x"008a1de5";
		wait for Clk_period;
		Addr <=  "00011101011100";
		Trees_din <= x"002a1de5";
		wait for Clk_period;
		Addr <=  "00011101011101";
		Trees_din <= x"06f77620";
		wait for Clk_period;
		Addr <=  "00011101011110";
		Trees_din <= x"0207bf10";
		wait for Clk_period;
		Addr <=  "00011101011111";
		Trees_din <= x"06f5f208";
		wait for Clk_period;
		Addr <=  "00011101100000";
		Trees_din <= x"09005804";
		wait for Clk_period;
		Addr <=  "00011101100001";
		Trees_din <= x"ff431de5";
		wait for Clk_period;
		Addr <=  "00011101100010";
		Trees_din <= x"004d1de5";
		wait for Clk_period;
		Addr <=  "00011101100011";
		Trees_din <= x"03fa1c04";
		wait for Clk_period;
		Addr <=  "00011101100100";
		Trees_din <= x"ffe71de5";
		wait for Clk_period;
		Addr <=  "00011101100101";
		Trees_din <= x"00a91de5";
		wait for Clk_period;
		Addr <=  "00011101100110";
		Trees_din <= x"04ff7608";
		wait for Clk_period;
		Addr <=  "00011101100111";
		Trees_din <= x"02094404";
		wait for Clk_period;
		Addr <=  "00011101101000";
		Trees_din <= x"00721de5";
		wait for Clk_period;
		Addr <=  "00011101101001";
		Trees_din <= x"00001de5";
		wait for Clk_period;
		Addr <=  "00011101101010";
		Trees_din <= x"15008204";
		wait for Clk_period;
		Addr <=  "00011101101011";
		Trees_din <= x"00161de5";
		wait for Clk_period;
		Addr <=  "00011101101100";
		Trees_din <= x"ff6f1de5";
		wait for Clk_period;
		Addr <=  "00011101101101";
		Trees_din <= x"0c002f04";
		wait for Clk_period;
		Addr <=  "00011101101110";
		Trees_din <= x"006d1de5";
		wait for Clk_period;
		Addr <=  "00011101101111";
		Trees_din <= x"1a00f108";
		wait for Clk_period;
		Addr <=  "00011101110000";
		Trees_din <= x"19008c04";
		wait for Clk_period;
		Addr <=  "00011101110001";
		Trees_din <= x"ffd01de5";
		wait for Clk_period;
		Addr <=  "00011101110010";
		Trees_din <= x"ff5c1de5";
		wait for Clk_period;
		Addr <=  "00011101110011";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00011101110100";
		Trees_din <= x"ffcd1de5";
		wait for Clk_period;
		Addr <=  "00011101110101";
		Trees_din <= x"00791de5";
		wait for Clk_period;
		Addr <=  "00011101110110";
		Trees_din <= x"1f000c04";
		wait for Clk_period;
		Addr <=  "00011101110111";
		Trees_din <= x"008a1de5";
		wait for Clk_period;
		Addr <=  "00011101111000";
		Trees_din <= x"ffd21de5";
		wait for Clk_period;
		Addr <=  "00011101111001";
		Trees_din <= x"00153250";
		wait for Clk_period;
		Addr <=  "00011101111010";
		Trees_din <= x"05011d38";
		wait for Clk_period;
		Addr <=  "00011101111011";
		Trees_din <= x"01fe261c";
		wait for Clk_period;
		Addr <=  "00011101111100";
		Trees_din <= x"05ff8110";
		wait for Clk_period;
		Addr <=  "00011101111101";
		Trees_din <= x"05fe9608";
		wait for Clk_period;
		Addr <=  "00011101111110";
		Trees_din <= x"08001b04";
		wait for Clk_period;
		Addr <=  "00011101111111";
		Trees_din <= x"ffc91ed9";
		wait for Clk_period;
		Addr <=  "00011110000000";
		Trees_din <= x"00491ed9";
		wait for Clk_period;
		Addr <=  "00011110000001";
		Trees_din <= x"09005204";
		wait for Clk_period;
		Addr <=  "00011110000010";
		Trees_din <= x"00231ed9";
		wait for Clk_period;
		Addr <=  "00011110000011";
		Trees_din <= x"ff711ed9";
		wait for Clk_period;
		Addr <=  "00011110000100";
		Trees_din <= x"16006504";
		wait for Clk_period;
		Addr <=  "00011110000101";
		Trees_din <= x"ffe61ed9";
		wait for Clk_period;
		Addr <=  "00011110000110";
		Trees_din <= x"03011204";
		wait for Clk_period;
		Addr <=  "00011110000111";
		Trees_din <= x"00c01ed9";
		wait for Clk_period;
		Addr <=  "00011110001000";
		Trees_din <= x"00051ed9";
		wait for Clk_period;
		Addr <=  "00011110001001";
		Trees_din <= x"05ffcd10";
		wait for Clk_period;
		Addr <=  "00011110001010";
		Trees_din <= x"0306c208";
		wait for Clk_period;
		Addr <=  "00011110001011";
		Trees_din <= x"1703f604";
		wait for Clk_period;
		Addr <=  "00011110001100";
		Trees_din <= x"00041ed9";
		wait for Clk_period;
		Addr <=  "00011110001101";
		Trees_din <= x"ffa31ed9";
		wait for Clk_period;
		Addr <=  "00011110001110";
		Trees_din <= x"1a00b404";
		wait for Clk_period;
		Addr <=  "00011110001111";
		Trees_din <= x"ffdc1ed9";
		wait for Clk_period;
		Addr <=  "00011110010000";
		Trees_din <= x"ff7c1ed9";
		wait for Clk_period;
		Addr <=  "00011110010001";
		Trees_din <= x"0d035308";
		wait for Clk_period;
		Addr <=  "00011110010010";
		Trees_din <= x"000ceb04";
		wait for Clk_period;
		Addr <=  "00011110010011";
		Trees_din <= x"ff5c1ed9";
		wait for Clk_period;
		Addr <=  "00011110010100";
		Trees_din <= x"ffcd1ed9";
		wait for Clk_period;
		Addr <=  "00011110010101";
		Trees_din <= x"003a1ed9";
		wait for Clk_period;
		Addr <=  "00011110010110";
		Trees_din <= x"0100bc10";
		wait for Clk_period;
		Addr <=  "00011110010111";
		Trees_din <= x"000fd30c";
		wait for Clk_period;
		Addr <=  "00011110011000";
		Trees_din <= x"06fe3308";
		wait for Clk_period;
		Addr <=  "00011110011001";
		Trees_din <= x"0bf98504";
		wait for Clk_period;
		Addr <=  "00011110011010";
		Trees_din <= x"ffeb1ed9";
		wait for Clk_period;
		Addr <=  "00011110011011";
		Trees_din <= x"ff571ed9";
		wait for Clk_period;
		Addr <=  "00011110011100";
		Trees_din <= x"fffb1ed9";
		wait for Clk_period;
		Addr <=  "00011110011101";
		Trees_din <= x"00061ed9";
		wait for Clk_period;
		Addr <=  "00011110011110";
		Trees_din <= x"07005804";
		wait for Clk_period;
		Addr <=  "00011110011111";
		Trees_din <= x"00101ed9";
		wait for Clk_period;
		Addr <=  "00011110100000";
		Trees_din <= x"00621ed9";
		wait for Clk_period;
		Addr <=  "00011110100001";
		Trees_din <= x"0bf9600c";
		wait for Clk_period;
		Addr <=  "00011110100010";
		Trees_din <= x"0f008308";
		wait for Clk_period;
		Addr <=  "00011110100011";
		Trees_din <= x"05f97204";
		wait for Clk_period;
		Addr <=  "00011110100100";
		Trees_din <= x"ff331ed9";
		wait for Clk_period;
		Addr <=  "00011110100101";
		Trees_din <= x"ffca1ed9";
		wait for Clk_period;
		Addr <=  "00011110100110";
		Trees_din <= x"00711ed9";
		wait for Clk_period;
		Addr <=  "00011110100111";
		Trees_din <= x"0e043e18";
		wait for Clk_period;
		Addr <=  "00011110101000";
		Trees_din <= x"13f83c08";
		wait for Clk_period;
		Addr <=  "00011110101001";
		Trees_din <= x"05fcdd04";
		wait for Clk_period;
		Addr <=  "00011110101010";
		Trees_din <= x"00281ed9";
		wait for Clk_period;
		Addr <=  "00011110101011";
		Trees_din <= x"ff6e1ed9";
		wait for Clk_period;
		Addr <=  "00011110101100";
		Trees_din <= x"010f0b08";
		wait for Clk_period;
		Addr <=  "00011110101101";
		Trees_din <= x"1900ab04";
		wait for Clk_period;
		Addr <=  "00011110101110";
		Trees_din <= x"007c1ed9";
		wait for Clk_period;
		Addr <=  "00011110101111";
		Trees_din <= x"00021ed9";
		wait for Clk_period;
		Addr <=  "00011110110000";
		Trees_din <= x"1d004a04";
		wait for Clk_period;
		Addr <=  "00011110110001";
		Trees_din <= x"003e1ed9";
		wait for Clk_period;
		Addr <=  "00011110110010";
		Trees_din <= x"ffc31ed9";
		wait for Clk_period;
		Addr <=  "00011110110011";
		Trees_din <= x"11043c04";
		wait for Clk_period;
		Addr <=  "00011110110100";
		Trees_din <= x"004b1ed9";
		wait for Clk_period;
		Addr <=  "00011110110101";
		Trees_din <= x"ff4f1ed9";
		wait for Clk_period;
		Addr <=  "00011110110110";
		Trees_din <= x"00229244";
		wait for Clk_period;
		Addr <=  "00011110110111";
		Trees_din <= x"09005e3c";
		wait for Clk_period;
		Addr <=  "00011110111000";
		Trees_din <= x"13f86f1c";
		wait for Clk_period;
		Addr <=  "00011110111001";
		Trees_din <= x"0efddb10";
		wait for Clk_period;
		Addr <=  "00011110111010";
		Trees_din <= x"13f7f008";
		wait for Clk_period;
		Addr <=  "00011110111011";
		Trees_din <= x"0b026f04";
		wait for Clk_period;
		Addr <=  "00011110111100";
		Trees_din <= x"00521f65";
		wait for Clk_period;
		Addr <=  "00011110111101";
		Trees_din <= x"ffee1f65";
		wait for Clk_period;
		Addr <=  "00011110111110";
		Trees_din <= x"1900a204";
		wait for Clk_period;
		Addr <=  "00011110111111";
		Trees_din <= x"ff5b1f65";
		wait for Clk_period;
		Addr <=  "00011111000000";
		Trees_din <= x"000a1f65";
		wait for Clk_period;
		Addr <=  "00011111000001";
		Trees_din <= x"09005708";
		wait for Clk_period;
		Addr <=  "00011111000010";
		Trees_din <= x"000c0a04";
		wait for Clk_period;
		Addr <=  "00011111000011";
		Trees_din <= x"00071f65";
		wait for Clk_period;
		Addr <=  "00011111000100";
		Trees_din <= x"00811f65";
		wait for Clk_period;
		Addr <=  "00011111000101";
		Trees_din <= x"ffb81f65";
		wait for Clk_period;
		Addr <=  "00011111000110";
		Trees_din <= x"13f8f710";
		wait for Clk_period;
		Addr <=  "00011111000111";
		Trees_din <= x"06f66008";
		wait for Clk_period;
		Addr <=  "00011111001000";
		Trees_din <= x"17039704";
		wait for Clk_period;
		Addr <=  "00011111001001";
		Trees_din <= x"00981f65";
		wait for Clk_period;
		Addr <=  "00011111001010";
		Trees_din <= x"ffa81f65";
		wait for Clk_period;
		Addr <=  "00011111001011";
		Trees_din <= x"19009e04";
		wait for Clk_period;
		Addr <=  "00011111001100";
		Trees_din <= x"ff991f65";
		wait for Clk_period;
		Addr <=  "00011111001101";
		Trees_din <= x"004f1f65";
		wait for Clk_period;
		Addr <=  "00011111001110";
		Trees_din <= x"1f000008";
		wait for Clk_period;
		Addr <=  "00011111001111";
		Trees_din <= x"04f47104";
		wait for Clk_period;
		Addr <=  "00011111010000";
		Trees_din <= x"004f1f65";
		wait for Clk_period;
		Addr <=  "00011111010001";
		Trees_din <= x"fff81f65";
		wait for Clk_period;
		Addr <=  "00011111010010";
		Trees_din <= x"07005304";
		wait for Clk_period;
		Addr <=  "00011111010011";
		Trees_din <= x"005a1f65";
		wait for Clk_period;
		Addr <=  "00011111010100";
		Trees_din <= x"fffc1f65";
		wait for Clk_period;
		Addr <=  "00011111010101";
		Trees_din <= x"01039c04";
		wait for Clk_period;
		Addr <=  "00011111010110";
		Trees_din <= x"ffd81f65";
		wait for Clk_period;
		Addr <=  "00011111010111";
		Trees_din <= x"008b1f65";
		wait for Clk_period;
		Addr <=  "00011111011000";
		Trees_din <= x"007e1f65";
		wait for Clk_period;
		Addr <=  "00011111011001";
		Trees_din <= x"00229248";
		wait for Clk_period;
		Addr <=  "00011111011010";
		Trees_din <= x"00fe7b08";
		wait for Clk_period;
		Addr <=  "00011111011011";
		Trees_din <= x"1f000004";
		wait for Clk_period;
		Addr <=  "00011111011100";
		Trees_din <= x"ff7e1ff9";
		wait for Clk_period;
		Addr <=  "00011111011101";
		Trees_din <= x"003f1ff9";
		wait for Clk_period;
		Addr <=  "00011111011110";
		Trees_din <= x"02071420";
		wait for Clk_period;
		Addr <=  "00011111011111";
		Trees_din <= x"06f3b410";
		wait for Clk_period;
		Addr <=  "00011111100000";
		Trees_din <= x"1603f708";
		wait for Clk_period;
		Addr <=  "00011111100001";
		Trees_din <= x"13015a04";
		wait for Clk_period;
		Addr <=  "00011111100010";
		Trees_din <= x"004f1ff9";
		wait for Clk_period;
		Addr <=  "00011111100011";
		Trees_din <= x"ffe51ff9";
		wait for Clk_period;
		Addr <=  "00011111100100";
		Trees_din <= x"06f2b704";
		wait for Clk_period;
		Addr <=  "00011111100101";
		Trees_din <= x"000f1ff9";
		wait for Clk_period;
		Addr <=  "00011111100110";
		Trees_din <= x"ff861ff9";
		wait for Clk_period;
		Addr <=  "00011111100111";
		Trees_din <= x"15009608";
		wait for Clk_period;
		Addr <=  "00011111101000";
		Trees_din <= x"0205dc04";
		wait for Clk_period;
		Addr <=  "00011111101001";
		Trees_din <= x"000f1ff9";
		wait for Clk_period;
		Addr <=  "00011111101010";
		Trees_din <= x"006a1ff9";
		wait for Clk_period;
		Addr <=  "00011111101011";
		Trees_din <= x"10f9ef04";
		wait for Clk_period;
		Addr <=  "00011111101100";
		Trees_din <= x"002d1ff9";
		wait for Clk_period;
		Addr <=  "00011111101101";
		Trees_din <= x"ffe81ff9";
		wait for Clk_period;
		Addr <=  "00011111101110";
		Trees_din <= x"0b04b810";
		wait for Clk_period;
		Addr <=  "00011111101111";
		Trees_din <= x"1b004208";
		wait for Clk_period;
		Addr <=  "00011111110000";
		Trees_din <= x"08001004";
		wait for Clk_period;
		Addr <=  "00011111110001";
		Trees_din <= x"00ac1ff9";
		wait for Clk_period;
		Addr <=  "00011111110010";
		Trees_din <= x"000e1ff9";
		wait for Clk_period;
		Addr <=  "00011111110011";
		Trees_din <= x"0c01c204";
		wait for Clk_period;
		Addr <=  "00011111110100";
		Trees_din <= x"00051ff9";
		wait for Clk_period;
		Addr <=  "00011111110101";
		Trees_din <= x"ff7b1ff9";
		wait for Clk_period;
		Addr <=  "00011111110110";
		Trees_din <= x"1b003f08";
		wait for Clk_period;
		Addr <=  "00011111110111";
		Trees_din <= x"2003ff04";
		wait for Clk_period;
		Addr <=  "00011111111000";
		Trees_din <= x"003f1ff9";
		wait for Clk_period;
		Addr <=  "00011111111001";
		Trees_din <= x"ff731ff9";
		wait for Clk_period;
		Addr <=  "00011111111010";
		Trees_din <= x"000f0704";
		wait for Clk_period;
		Addr <=  "00011111111011";
		Trees_din <= x"ffa31ff9";
		wait for Clk_period;
		Addr <=  "00011111111100";
		Trees_din <= x"007c1ff9";
		wait for Clk_period;
		Addr <=  "00011111111101";
		Trees_din <= x"00791ff9";
		wait for Clk_period;
		Addr <=  "00011111111110";
		Trees_din <= x"0003aa34";
		wait for Clk_period;
		Addr <=  "00011111111111";
		Trees_din <= x"1b003d18";
		wait for Clk_period;
		Addr <=  "00100000000000";
		Trees_din <= x"08022f0c";
		wait for Clk_period;
		Addr <=  "00100000000001";
		Trees_din <= x"10f72e04";
		wait for Clk_period;
		Addr <=  "00100000000010";
		Trees_din <= x"003a2115";
		wait for Clk_period;
		Addr <=  "00100000000011";
		Trees_din <= x"02fba504";
		wait for Clk_period;
		Addr <=  "00100000000100";
		Trees_din <= x"000a2115";
		wait for Clk_period;
		Addr <=  "00100000000101";
		Trees_din <= x"ff702115";
		wait for Clk_period;
		Addr <=  "00100000000110";
		Trees_din <= x"0afde308";
		wait for Clk_period;
		Addr <=  "00100000000111";
		Trees_din <= x"13ffe604";
		wait for Clk_period;
		Addr <=  "00100000001000";
		Trees_din <= x"00992115";
		wait for Clk_period;
		Addr <=  "00100000001001";
		Trees_din <= x"00032115";
		wait for Clk_period;
		Addr <=  "00100000001010";
		Trees_din <= x"ff8d2115";
		wait for Clk_period;
		Addr <=  "00100000001011";
		Trees_din <= x"07005814";
		wait for Clk_period;
		Addr <=  "00100000001100";
		Trees_din <= x"08001a04";
		wait for Clk_period;
		Addr <=  "00100000001101";
		Trees_din <= x"ffa42115";
		wait for Clk_period;
		Addr <=  "00100000001110";
		Trees_din <= x"07005508";
		wait for Clk_period;
		Addr <=  "00100000001111";
		Trees_din <= x"01fb9304";
		wait for Clk_period;
		Addr <=  "00100000010000";
		Trees_din <= x"00592115";
		wait for Clk_period;
		Addr <=  "00100000010001";
		Trees_din <= x"ffb62115";
		wait for Clk_period;
		Addr <=  "00100000010010";
		Trees_din <= x"1b003f04";
		wait for Clk_period;
		Addr <=  "00100000010011";
		Trees_din <= x"00c82115";
		wait for Clk_period;
		Addr <=  "00100000010100";
		Trees_din <= x"003b2115";
		wait for Clk_period;
		Addr <=  "00100000010101";
		Trees_din <= x"15009c04";
		wait for Clk_period;
		Addr <=  "00100000010110";
		Trees_din <= x"ff862115";
		wait for Clk_period;
		Addr <=  "00100000010111";
		Trees_din <= x"00272115";
		wait for Clk_period;
		Addr <=  "00100000011000";
		Trees_din <= x"02fdcd1c";
		wait for Clk_period;
		Addr <=  "00100000011001";
		Trees_din <= x"01082a10";
		wait for Clk_period;
		Addr <=  "00100000011010";
		Trees_din <= x"05fe640c";
		wait for Clk_period;
		Addr <=  "00100000011011";
		Trees_din <= x"0bf97c04";
		wait for Clk_period;
		Addr <=  "00100000011100";
		Trees_din <= x"00142115";
		wait for Clk_period;
		Addr <=  "00100000011101";
		Trees_din <= x"1600af04";
		wait for Clk_period;
		Addr <=  "00100000011110";
		Trees_din <= x"00202115";
		wait for Clk_period;
		Addr <=  "00100000011111";
		Trees_din <= x"00982115";
		wait for Clk_period;
		Addr <=  "00100000100000";
		Trees_din <= x"fffd2115";
		wait for Clk_period;
		Addr <=  "00100000100001";
		Trees_din <= x"09005808";
		wait for Clk_period;
		Addr <=  "00100000100010";
		Trees_din <= x"02fd8004";
		wait for Clk_period;
		Addr <=  "00100000100011";
		Trees_din <= x"ff9f2115";
		wait for Clk_period;
		Addr <=  "00100000100100";
		Trees_din <= x"00262115";
		wait for Clk_period;
		Addr <=  "00100000100101";
		Trees_din <= x"005f2115";
		wait for Clk_period;
		Addr <=  "00100000100110";
		Trees_din <= x"08000f20";
		wait for Clk_period;
		Addr <=  "00100000100111";
		Trees_din <= x"1200c310";
		wait for Clk_period;
		Addr <=  "00100000101000";
		Trees_din <= x"11fef808";
		wait for Clk_period;
		Addr <=  "00100000101001";
		Trees_din <= x"0c018304";
		wait for Clk_period;
		Addr <=  "00100000101010";
		Trees_din <= x"006d2115";
		wait for Clk_period;
		Addr <=  "00100000101011";
		Trees_din <= x"ff972115";
		wait for Clk_period;
		Addr <=  "00100000101100";
		Trees_din <= x"0d00a704";
		wait for Clk_period;
		Addr <=  "00100000101101";
		Trees_din <= x"000a2115";
		wait for Clk_period;
		Addr <=  "00100000101110";
		Trees_din <= x"00a32115";
		wait for Clk_period;
		Addr <=  "00100000101111";
		Trees_din <= x"07005608";
		wait for Clk_period;
		Addr <=  "00100000110000";
		Trees_din <= x"010fd304";
		wait for Clk_period;
		Addr <=  "00100000110001";
		Trees_din <= x"00982115";
		wait for Clk_period;
		Addr <=  "00100000110010";
		Trees_din <= x"ffc52115";
		wait for Clk_period;
		Addr <=  "00100000110011";
		Trees_din <= x"1a00b804";
		wait for Clk_period;
		Addr <=  "00100000110100";
		Trees_din <= x"00122115";
		wait for Clk_period;
		Addr <=  "00100000110101";
		Trees_din <= x"ff862115";
		wait for Clk_period;
		Addr <=  "00100000110110";
		Trees_din <= x"18004810";
		wait for Clk_period;
		Addr <=  "00100000110111";
		Trees_din <= x"15009208";
		wait for Clk_period;
		Addr <=  "00100000111000";
		Trees_din <= x"04fc8204";
		wait for Clk_period;
		Addr <=  "00100000111001";
		Trees_din <= x"000c2115";
		wait for Clk_period;
		Addr <=  "00100000111010";
		Trees_din <= x"00712115";
		wait for Clk_period;
		Addr <=  "00100000111011";
		Trees_din <= x"0d02e504";
		wait for Clk_period;
		Addr <=  "00100000111100";
		Trees_din <= x"000b2115";
		wait for Clk_period;
		Addr <=  "00100000111101";
		Trees_din <= x"ffde2115";
		wait for Clk_period;
		Addr <=  "00100000111110";
		Trees_din <= x"00108808";
		wait for Clk_period;
		Addr <=  "00100000111111";
		Trees_din <= x"05fbfd04";
		wait for Clk_period;
		Addr <=  "00100001000000";
		Trees_din <= x"ff9f2115";
		wait for Clk_period;
		Addr <=  "00100001000001";
		Trees_din <= x"00082115";
		wait for Clk_period;
		Addr <=  "00100001000010";
		Trees_din <= x"1b003f04";
		wait for Clk_period;
		Addr <=  "00100001000011";
		Trees_din <= x"ffc22115";
		wait for Clk_period;
		Addr <=  "00100001000100";
		Trees_din <= x"002a2115";
		wait for Clk_period;
		Addr <=  "00100001000101";
		Trees_din <= x"00229230";
		wait for Clk_period;
		Addr <=  "00100001000110";
		Trees_din <= x"09005e28";
		wait for Clk_period;
		Addr <=  "00100001000111";
		Trees_din <= x"09005d20";
		wait for Clk_period;
		Addr <=  "00100001001000";
		Trees_din <= x"13f86f10";
		wait for Clk_period;
		Addr <=  "00100001001001";
		Trees_din <= x"1400c508";
		wait for Clk_period;
		Addr <=  "00100001001010";
		Trees_din <= x"0f001304";
		wait for Clk_period;
		Addr <=  "00100001001011";
		Trees_din <= x"ffd72179";
		wait for Clk_period;
		Addr <=  "00100001001100";
		Trees_din <= x"00552179";
		wait for Clk_period;
		Addr <=  "00100001001101";
		Trees_din <= x"18003e04";
		wait for Clk_period;
		Addr <=  "00100001001110";
		Trees_din <= x"00332179";
		wait for Clk_period;
		Addr <=  "00100001001111";
		Trees_din <= x"ff622179";
		wait for Clk_period;
		Addr <=  "00100001010000";
		Trees_din <= x"13f8f708";
		wait for Clk_period;
		Addr <=  "00100001010001";
		Trees_din <= x"06f66004";
		wait for Clk_period;
		Addr <=  "00100001010010";
		Trees_din <= x"00632179";
		wait for Clk_period;
		Addr <=  "00100001010011";
		Trees_din <= x"ffd52179";
		wait for Clk_period;
		Addr <=  "00100001010100";
		Trees_din <= x"07005b04";
		wait for Clk_period;
		Addr <=  "00100001010101";
		Trees_din <= x"00042179";
		wait for Clk_period;
		Addr <=  "00100001010110";
		Trees_din <= x"ffe12179";
		wait for Clk_period;
		Addr <=  "00100001010111";
		Trees_din <= x"1a00bc04";
		wait for Clk_period;
		Addr <=  "00100001011000";
		Trees_din <= x"00002179";
		wait for Clk_period;
		Addr <=  "00100001011001";
		Trees_din <= x"ff612179";
		wait for Clk_period;
		Addr <=  "00100001011010";
		Trees_din <= x"01039c04";
		wait for Clk_period;
		Addr <=  "00100001011011";
		Trees_din <= x"ffdd2179";
		wait for Clk_period;
		Addr <=  "00100001011100";
		Trees_din <= x"00802179";
		wait for Clk_period;
		Addr <=  "00100001011101";
		Trees_din <= x"00712179";
		wait for Clk_period;
		Addr <=  "00100001011110";
		Trees_din <= x"00153240";
		wait for Clk_period;
		Addr <=  "00100001011111";
		Trees_din <= x"0bf90c1c";
		wait for Clk_period;
		Addr <=  "00100001100000";
		Trees_din <= x"09005008";
		wait for Clk_period;
		Addr <=  "00100001100001";
		Trees_din <= x"07005204";
		wait for Clk_period;
		Addr <=  "00100001100010";
		Trees_din <= x"00222255";
		wait for Clk_period;
		Addr <=  "00100001100011";
		Trees_din <= x"ff672255";
		wait for Clk_period;
		Addr <=  "00100001100100";
		Trees_din <= x"000bca08";
		wait for Clk_period;
		Addr <=  "00100001100101";
		Trees_din <= x"1003e904";
		wait for Clk_period;
		Addr <=  "00100001100110";
		Trees_din <= x"00682255";
		wait for Clk_period;
		Addr <=  "00100001100111";
		Trees_din <= x"ffa22255";
		wait for Clk_period;
		Addr <=  "00100001101000";
		Trees_din <= x"0f02d608";
		wait for Clk_period;
		Addr <=  "00100001101001";
		Trees_din <= x"1c002d04";
		wait for Clk_period;
		Addr <=  "00100001101010";
		Trees_din <= x"001d2255";
		wait for Clk_period;
		Addr <=  "00100001101011";
		Trees_din <= x"00b82255";
		wait for Clk_period;
		Addr <=  "00100001101100";
		Trees_din <= x"ffbd2255";
		wait for Clk_period;
		Addr <=  "00100001101101";
		Trees_din <= x"03f23604";
		wait for Clk_period;
		Addr <=  "00100001101110";
		Trees_din <= x"00712255";
		wait for Clk_period;
		Addr <=  "00100001101111";
		Trees_din <= x"02094410";
		wait for Clk_period;
		Addr <=  "00100001110000";
		Trees_din <= x"06f63b08";
		wait for Clk_period;
		Addr <=  "00100001110001";
		Trees_din <= x"05fede04";
		wait for Clk_period;
		Addr <=  "00100001110010";
		Trees_din <= x"00142255";
		wait for Clk_period;
		Addr <=  "00100001110011";
		Trees_din <= x"ff982255";
		wait for Clk_period;
		Addr <=  "00100001110100";
		Trees_din <= x"0d02e504";
		wait for Clk_period;
		Addr <=  "00100001110101";
		Trees_din <= x"00042255";
		wait for Clk_period;
		Addr <=  "00100001110110";
		Trees_din <= x"ffcd2255";
		wait for Clk_period;
		Addr <=  "00100001110111";
		Trees_din <= x"08008508";
		wait for Clk_period;
		Addr <=  "00100001111000";
		Trees_din <= x"1e006d04";
		wait for Clk_period;
		Addr <=  "00100001111001";
		Trees_din <= x"00952255";
		wait for Clk_period;
		Addr <=  "00100001111010";
		Trees_din <= x"ffc32255";
		wait for Clk_period;
		Addr <=  "00100001111011";
		Trees_din <= x"0bfa4104";
		wait for Clk_period;
		Addr <=  "00100001111100";
		Trees_din <= x"ff5f2255";
		wait for Clk_period;
		Addr <=  "00100001111101";
		Trees_din <= x"ffd32255";
		wait for Clk_period;
		Addr <=  "00100001111110";
		Trees_din <= x"0bf9600c";
		wait for Clk_period;
		Addr <=  "00100001111111";
		Trees_din <= x"0f008308";
		wait for Clk_period;
		Addr <=  "00100010000000";
		Trees_din <= x"07005804";
		wait for Clk_period;
		Addr <=  "00100010000001";
		Trees_din <= x"ff5c2255";
		wait for Clk_period;
		Addr <=  "00100010000010";
		Trees_din <= x"ffdf2255";
		wait for Clk_period;
		Addr <=  "00100010000011";
		Trees_din <= x"00672255";
		wait for Clk_period;
		Addr <=  "00100010000100";
		Trees_din <= x"0f007f08";
		wait for Clk_period;
		Addr <=  "00100010000101";
		Trees_din <= x"05fe5c04";
		wait for Clk_period;
		Addr <=  "00100010000110";
		Trees_din <= x"007f2255";
		wait for Clk_period;
		Addr <=  "00100010000111";
		Trees_din <= x"00132255";
		wait for Clk_period;
		Addr <=  "00100010001000";
		Trees_din <= x"1c00310c";
		wait for Clk_period;
		Addr <=  "00100010001001";
		Trees_din <= x"0f03ba08";
		wait for Clk_period;
		Addr <=  "00100010001010";
		Trees_din <= x"16037404";
		wait for Clk_period;
		Addr <=  "00100010001011";
		Trees_din <= x"006d2255";
		wait for Clk_period;
		Addr <=  "00100010001100";
		Trees_din <= x"ffc42255";
		wait for Clk_period;
		Addr <=  "00100010001101";
		Trees_din <= x"ff492255";
		wait for Clk_period;
		Addr <=  "00100010001110";
		Trees_din <= x"03f2cc08";
		wait for Clk_period;
		Addr <=  "00100010001111";
		Trees_din <= x"17000004";
		wait for Clk_period;
		Addr <=  "00100010010000";
		Trees_din <= x"00492255";
		wait for Clk_period;
		Addr <=  "00100010010001";
		Trees_din <= x"ffa62255";
		wait for Clk_period;
		Addr <=  "00100010010010";
		Trees_din <= x"0c035e04";
		wait for Clk_period;
		Addr <=  "00100010010011";
		Trees_din <= x"007b2255";
		wait for Clk_period;
		Addr <=  "00100010010100";
		Trees_din <= x"ffe72255";
		wait for Clk_period;
		Addr <=  "00100010010101";
		Trees_din <= x"0007905c";
		wait for Clk_period;
		Addr <=  "00100010010110";
		Trees_din <= x"13ffd534";
		wait for Clk_period;
		Addr <=  "00100010010111";
		Trees_din <= x"1102881c";
		wait for Clk_period;
		Addr <=  "00100010011000";
		Trees_din <= x"17018e0c";
		wait for Clk_period;
		Addr <=  "00100010011001";
		Trees_din <= x"0e02bd08";
		wait for Clk_period;
		Addr <=  "00100010011010";
		Trees_din <= x"00072f04";
		wait for Clk_period;
		Addr <=  "00100010011011";
		Trees_din <= x"ff8423c9";
		wait for Clk_period;
		Addr <=  "00100010011100";
		Trees_din <= x"002123c9";
		wait for Clk_period;
		Addr <=  "00100010011101";
		Trees_din <= x"004223c9";
		wait for Clk_period;
		Addr <=  "00100010011110";
		Trees_din <= x"07005808";
		wait for Clk_period;
		Addr <=  "00100010011111";
		Trees_din <= x"01fec704";
		wait for Clk_period;
		Addr <=  "00100010100000";
		Trees_din <= x"001423c9";
		wait for Clk_period;
		Addr <=  "00100010100001";
		Trees_din <= x"ff7d23c9";
		wait for Clk_period;
		Addr <=  "00100010100010";
		Trees_din <= x"0d01fd04";
		wait for Clk_period;
		Addr <=  "00100010100011";
		Trees_din <= x"fff723c9";
		wait for Clk_period;
		Addr <=  "00100010100100";
		Trees_din <= x"00a223c9";
		wait for Clk_period;
		Addr <=  "00100010100101";
		Trees_din <= x"17005c10";
		wait for Clk_period;
		Addr <=  "00100010100110";
		Trees_din <= x"09005408";
		wait for Clk_period;
		Addr <=  "00100010100111";
		Trees_din <= x"09005004";
		wait for Clk_period;
		Addr <=  "00100010101000";
		Trees_din <= x"003a23c9";
		wait for Clk_period;
		Addr <=  "00100010101001";
		Trees_din <= x"00d923c9";
		wait for Clk_period;
		Addr <=  "00100010101010";
		Trees_din <= x"0403b004";
		wait for Clk_period;
		Addr <=  "00100010101011";
		Trees_din <= x"ff9123c9";
		wait for Clk_period;
		Addr <=  "00100010101100";
		Trees_din <= x"006323c9";
		wait for Clk_period;
		Addr <=  "00100010101101";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00100010101110";
		Trees_din <= x"ff7723c9";
		wait for Clk_period;
		Addr <=  "00100010101111";
		Trees_din <= x"000523c9";
		wait for Clk_period;
		Addr <=  "00100010110000";
		Trees_din <= x"07005618";
		wait for Clk_period;
		Addr <=  "00100010110001";
		Trees_din <= x"0bfa3808";
		wait for Clk_period;
		Addr <=  "00100010110010";
		Trees_din <= x"11023204";
		wait for Clk_period;
		Addr <=  "00100010110011";
		Trees_din <= x"00ab23c9";
		wait for Clk_period;
		Addr <=  "00100010110100";
		Trees_din <= x"002323c9";
		wait for Clk_period;
		Addr <=  "00100010110101";
		Trees_din <= x"0d017008";
		wait for Clk_period;
		Addr <=  "00100010110110";
		Trees_din <= x"09005104";
		wait for Clk_period;
		Addr <=  "00100010110111";
		Trees_din <= x"ffe923c9";
		wait for Clk_period;
		Addr <=  "00100010111000";
		Trees_din <= x"008623c9";
		wait for Clk_period;
		Addr <=  "00100010111001";
		Trees_din <= x"17000204";
		wait for Clk_period;
		Addr <=  "00100010111010";
		Trees_din <= x"002623c9";
		wait for Clk_period;
		Addr <=  "00100010111011";
		Trees_din <= x"ffa223c9";
		wait for Clk_period;
		Addr <=  "00100010111100";
		Trees_din <= x"05fd1d04";
		wait for Clk_period;
		Addr <=  "00100010111101";
		Trees_din <= x"ff7723c9";
		wait for Clk_period;
		Addr <=  "00100010111110";
		Trees_din <= x"03ff7d04";
		wait for Clk_period;
		Addr <=  "00100010111111";
		Trees_din <= x"ffc323c9";
		wait for Clk_period;
		Addr <=  "00100011000000";
		Trees_din <= x"0204d704";
		wait for Clk_period;
		Addr <=  "00100011000001";
		Trees_din <= x"001423c9";
		wait for Clk_period;
		Addr <=  "00100011000010";
		Trees_din <= x"009023c9";
		wait for Clk_period;
		Addr <=  "00100011000011";
		Trees_din <= x"04ff5740";
		wait for Clk_period;
		Addr <=  "00100011000100";
		Trees_din <= x"0102bb20";
		wait for Clk_period;
		Addr <=  "00100011000101";
		Trees_din <= x"13fa6410";
		wait for Clk_period;
		Addr <=  "00100011000110";
		Trees_din <= x"1c003108";
		wait for Clk_period;
		Addr <=  "00100011000111";
		Trees_din <= x"05007904";
		wait for Clk_period;
		Addr <=  "00100011001000";
		Trees_din <= x"005b23c9";
		wait for Clk_period;
		Addr <=  "00100011001001";
		Trees_din <= x"ffdf23c9";
		wait for Clk_period;
		Addr <=  "00100011001010";
		Trees_din <= x"00138a04";
		wait for Clk_period;
		Addr <=  "00100011001011";
		Trees_din <= x"ff8123c9";
		wait for Clk_period;
		Addr <=  "00100011001100";
		Trees_din <= x"001e23c9";
		wait for Clk_period;
		Addr <=  "00100011001101";
		Trees_din <= x"05fff708";
		wait for Clk_period;
		Addr <=  "00100011001110";
		Trees_din <= x"07005504";
		wait for Clk_period;
		Addr <=  "00100011001111";
		Trees_din <= x"001423c9";
		wait for Clk_period;
		Addr <=  "00100011010000";
		Trees_din <= x"008623c9";
		wait for Clk_period;
		Addr <=  "00100011010001";
		Trees_din <= x"0bfa8d04";
		wait for Clk_period;
		Addr <=  "00100011010010";
		Trees_din <= x"005923c9";
		wait for Clk_period;
		Addr <=  "00100011010011";
		Trees_din <= x"ffab23c9";
		wait for Clk_period;
		Addr <=  "00100011010100";
		Trees_din <= x"08001710";
		wait for Clk_period;
		Addr <=  "00100011010101";
		Trees_din <= x"06f96108";
		wait for Clk_period;
		Addr <=  "00100011010110";
		Trees_din <= x"01139004";
		wait for Clk_period;
		Addr <=  "00100011010111";
		Trees_din <= x"005723c9";
		wait for Clk_period;
		Addr <=  "00100011011000";
		Trees_din <= x"ffab23c9";
		wait for Clk_period;
		Addr <=  "00100011011001";
		Trees_din <= x"05fa9804";
		wait for Clk_period;
		Addr <=  "00100011011010";
		Trees_din <= x"ff5823c9";
		wait for Clk_period;
		Addr <=  "00100011011011";
		Trees_din <= x"005323c9";
		wait for Clk_period;
		Addr <=  "00100011011100";
		Trees_din <= x"03fb7408";
		wait for Clk_period;
		Addr <=  "00100011011101";
		Trees_din <= x"0bfad104";
		wait for Clk_period;
		Addr <=  "00100011011110";
		Trees_din <= x"ffdd23c9";
		wait for Clk_period;
		Addr <=  "00100011011111";
		Trees_din <= x"000a23c9";
		wait for Clk_period;
		Addr <=  "00100011100000";
		Trees_din <= x"1402a204";
		wait for Clk_period;
		Addr <=  "00100011100001";
		Trees_din <= x"ffa923c9";
		wait for Clk_period;
		Addr <=  "00100011100010";
		Trees_din <= x"001c23c9";
		wait for Clk_period;
		Addr <=  "00100011100011";
		Trees_din <= x"07005a10";
		wait for Clk_period;
		Addr <=  "00100011100100";
		Trees_din <= x"08000b04";
		wait for Clk_period;
		Addr <=  "00100011100101";
		Trees_din <= x"ff6723c9";
		wait for Clk_period;
		Addr <=  "00100011100110";
		Trees_din <= x"10f90b04";
		wait for Clk_period;
		Addr <=  "00100011100111";
		Trees_din <= x"009823c9";
		wait for Clk_period;
		Addr <=  "00100011101000";
		Trees_din <= x"010b8f04";
		wait for Clk_period;
		Addr <=  "00100011101001";
		Trees_din <= x"002623c9";
		wait for Clk_period;
		Addr <=  "00100011101010";
		Trees_din <= x"ff9523c9";
		wait for Clk_period;
		Addr <=  "00100011101011";
		Trees_din <= x"1c004108";
		wait for Clk_period;
		Addr <=  "00100011101100";
		Trees_din <= x"1b003304";
		wait for Clk_period;
		Addr <=  "00100011101101";
		Trees_din <= x"ffcf23c9";
		wait for Clk_period;
		Addr <=  "00100011101110";
		Trees_din <= x"00b823c9";
		wait for Clk_period;
		Addr <=  "00100011101111";
		Trees_din <= x"0c01c204";
		wait for Clk_period;
		Addr <=  "00100011110000";
		Trees_din <= x"ff8f23c9";
		wait for Clk_period;
		Addr <=  "00100011110001";
		Trees_din <= x"004823c9";
		wait for Clk_period;
		Addr <=  "00100011110010";
		Trees_din <= x"000f6f6c";
		wait for Clk_period;
		Addr <=  "00100011110011";
		Trees_din <= x"19008330";
		wait for Clk_period;
		Addr <=  "00100011110100";
		Trees_din <= x"05fc1218";
		wait for Clk_period;
		Addr <=  "00100011110101";
		Trees_din <= x"0a044c10";
		wait for Clk_period;
		Addr <=  "00100011110110";
		Trees_din <= x"08002d08";
		wait for Clk_period;
		Addr <=  "00100011110111";
		Trees_din <= x"06f37f04";
		wait for Clk_period;
		Addr <=  "00100011111000";
		Trees_din <= x"0053253d";
		wait for Clk_period;
		Addr <=  "00100011111001";
		Trees_din <= x"ffa7253d";
		wait for Clk_period;
		Addr <=  "00100011111010";
		Trees_din <= x"04007b04";
		wait for Clk_period;
		Addr <=  "00100011111011";
		Trees_din <= x"ff61253d";
		wait for Clk_period;
		Addr <=  "00100011111100";
		Trees_din <= x"ffca253d";
		wait for Clk_period;
		Addr <=  "00100011111101";
		Trees_din <= x"10fade04";
		wait for Clk_period;
		Addr <=  "00100011111110";
		Trees_din <= x"0085253d";
		wait for Clk_period;
		Addr <=  "00100011111111";
		Trees_din <= x"ffe4253d";
		wait for Clk_period;
		Addr <=  "00100100000000";
		Trees_din <= x"01077d10";
		wait for Clk_period;
		Addr <=  "00100100000001";
		Trees_din <= x"02ff9d08";
		wait for Clk_period;
		Addr <=  "00100100000010";
		Trees_din <= x"11005c04";
		wait for Clk_period;
		Addr <=  "00100100000011";
		Trees_din <= x"005b253d";
		wait for Clk_period;
		Addr <=  "00100100000100";
		Trees_din <= x"0017253d";
		wait for Clk_period;
		Addr <=  "00100100000101";
		Trees_din <= x"11028804";
		wait for Clk_period;
		Addr <=  "00100100000110";
		Trees_din <= x"ff80253d";
		wait for Clk_period;
		Addr <=  "00100100000111";
		Trees_din <= x"000c253d";
		wait for Clk_period;
		Addr <=  "00100100001000";
		Trees_din <= x"06f3ec04";
		wait for Clk_period;
		Addr <=  "00100100001001";
		Trees_din <= x"ffe8253d";
		wait for Clk_period;
		Addr <=  "00100100001010";
		Trees_din <= x"00a0253d";
		wait for Clk_period;
		Addr <=  "00100100001011";
		Trees_din <= x"1c003d20";
		wait for Clk_period;
		Addr <=  "00100100001100";
		Trees_din <= x"000e9010";
		wait for Clk_period;
		Addr <=  "00100100001101";
		Trees_din <= x"1004a908";
		wait for Clk_period;
		Addr <=  "00100100001110";
		Trees_din <= x"1b002f04";
		wait for Clk_period;
		Addr <=  "00100100001111";
		Trees_din <= x"ffd4253d";
		wait for Clk_period;
		Addr <=  "00100100010000";
		Trees_din <= x"001d253d";
		wait for Clk_period;
		Addr <=  "00100100010001";
		Trees_din <= x"08002104";
		wait for Clk_period;
		Addr <=  "00100100010010";
		Trees_din <= x"0048253d";
		wait for Clk_period;
		Addr <=  "00100100010011";
		Trees_din <= x"ffcb253d";
		wait for Clk_period;
		Addr <=  "00100100010100";
		Trees_din <= x"16002d08";
		wait for Clk_period;
		Addr <=  "00100100010101";
		Trees_din <= x"07005a04";
		wait for Clk_period;
		Addr <=  "00100100010110";
		Trees_din <= x"007a253d";
		wait for Clk_period;
		Addr <=  "00100100010111";
		Trees_din <= x"ffd8253d";
		wait for Clk_period;
		Addr <=  "00100100011000";
		Trees_din <= x"06f1ee04";
		wait for Clk_period;
		Addr <=  "00100100011001";
		Trees_din <= x"006b253d";
		wait for Clk_period;
		Addr <=  "00100100011010";
		Trees_din <= x"ff85253d";
		wait for Clk_period;
		Addr <=  "00100100011011";
		Trees_din <= x"010b320c";
		wait for Clk_period;
		Addr <=  "00100100011100";
		Trees_din <= x"0d011d04";
		wait for Clk_period;
		Addr <=  "00100100011101";
		Trees_din <= x"ff6a253d";
		wait for Clk_period;
		Addr <=  "00100100011110";
		Trees_din <= x"1e007604";
		wait for Clk_period;
		Addr <=  "00100100011111";
		Trees_din <= x"ffac253d";
		wait for Clk_period;
		Addr <=  "00100100100000";
		Trees_din <= x"0062253d";
		wait for Clk_period;
		Addr <=  "00100100100001";
		Trees_din <= x"010fd308";
		wait for Clk_period;
		Addr <=  "00100100100010";
		Trees_din <= x"04fe3404";
		wait for Clk_period;
		Addr <=  "00100100100011";
		Trees_din <= x"00f0253d";
		wait for Clk_period;
		Addr <=  "00100100100100";
		Trees_din <= x"0008253d";
		wait for Clk_period;
		Addr <=  "00100100100101";
		Trees_din <= x"1b004604";
		wait for Clk_period;
		Addr <=  "00100100100110";
		Trees_din <= x"ffa8253d";
		wait for Clk_period;
		Addr <=  "00100100100111";
		Trees_din <= x"005b253d";
		wait for Clk_period;
		Addr <=  "00100100101000";
		Trees_din <= x"0afb0124";
		wait for Clk_period;
		Addr <=  "00100100101001";
		Trees_din <= x"11009a04";
		wait for Clk_period;
		Addr <=  "00100100101010";
		Trees_din <= x"008a253d";
		wait for Clk_period;
		Addr <=  "00100100101011";
		Trees_din <= x"17000310";
		wait for Clk_period;
		Addr <=  "00100100101100";
		Trees_din <= x"07005808";
		wait for Clk_period;
		Addr <=  "00100100101101";
		Trees_din <= x"07005504";
		wait for Clk_period;
		Addr <=  "00100100101110";
		Trees_din <= x"ffd9253d";
		wait for Clk_period;
		Addr <=  "00100100101111";
		Trees_din <= x"ff19253d";
		wait for Clk_period;
		Addr <=  "00100100110000";
		Trees_din <= x"0b043804";
		wait for Clk_period;
		Addr <=  "00100100110001";
		Trees_din <= x"0078253d";
		wait for Clk_period;
		Addr <=  "00100100110010";
		Trees_din <= x"ff9d253d";
		wait for Clk_period;
		Addr <=  "00100100110011";
		Trees_din <= x"00119208";
		wait for Clk_period;
		Addr <=  "00100100110100";
		Trees_din <= x"10043304";
		wait for Clk_period;
		Addr <=  "00100100110101";
		Trees_din <= x"ff7a253d";
		wait for Clk_period;
		Addr <=  "00100100110110";
		Trees_din <= x"0045253d";
		wait for Clk_period;
		Addr <=  "00100100110111";
		Trees_din <= x"05f82b04";
		wait for Clk_period;
		Addr <=  "00100100111000";
		Trees_din <= x"ffbb253d";
		wait for Clk_period;
		Addr <=  "00100100111001";
		Trees_din <= x"0045253d";
		wait for Clk_period;
		Addr <=  "00100100111010";
		Trees_din <= x"0afb260c";
		wait for Clk_period;
		Addr <=  "00100100111011";
		Trees_din <= x"0c00ed08";
		wait for Clk_period;
		Addr <=  "00100100111100";
		Trees_din <= x"1603e304";
		wait for Clk_period;
		Addr <=  "00100100111101";
		Trees_din <= x"ff62253d";
		wait for Clk_period;
		Addr <=  "00100100111110";
		Trees_din <= x"0052253d";
		wait for Clk_period;
		Addr <=  "00100100111111";
		Trees_din <= x"00ac253d";
		wait for Clk_period;
		Addr <=  "00100101000000";
		Trees_din <= x"09005a10";
		wait for Clk_period;
		Addr <=  "00100101000001";
		Trees_din <= x"0c036408";
		wait for Clk_period;
		Addr <=  "00100101000010";
		Trees_din <= x"0203ea04";
		wait for Clk_period;
		Addr <=  "00100101000011";
		Trees_din <= x"004c253d";
		wait for Clk_period;
		Addr <=  "00100101000100";
		Trees_din <= x"0006253d";
		wait for Clk_period;
		Addr <=  "00100101000101";
		Trees_din <= x"1e008104";
		wait for Clk_period;
		Addr <=  "00100101000110";
		Trees_din <= x"ffbe253d";
		wait for Clk_period;
		Addr <=  "00100101000111";
		Trees_din <= x"0073253d";
		wait for Clk_period;
		Addr <=  "00100101001000";
		Trees_din <= x"11028708";
		wait for Clk_period;
		Addr <=  "00100101001001";
		Trees_din <= x"03f52404";
		wait for Clk_period;
		Addr <=  "00100101001010";
		Trees_din <= x"ffa0253d";
		wait for Clk_period;
		Addr <=  "00100101001011";
		Trees_din <= x"0054253d";
		wait for Clk_period;
		Addr <=  "00100101001100";
		Trees_din <= x"06f69e04";
		wait for Clk_period;
		Addr <=  "00100101001101";
		Trees_din <= x"ff41253d";
		wait for Clk_period;
		Addr <=  "00100101001110";
		Trees_din <= x"0003253d";
		wait for Clk_period;
		Addr <=  "00100101001111";
		Trees_din <= x"02071458";
		wait for Clk_period;
		Addr <=  "00100101010000";
		Trees_din <= x"04f6cb24";
		wait for Clk_period;
		Addr <=  "00100101010001";
		Trees_din <= x"0afaf60c";
		wait for Clk_period;
		Addr <=  "00100101010010";
		Trees_din <= x"1b003604";
		wait for Clk_period;
		Addr <=  "00100101010011";
		Trees_din <= x"ff5d2691";
		wait for Clk_period;
		Addr <=  "00100101010100";
		Trees_din <= x"0011ff04";
		wait for Clk_period;
		Addr <=  "00100101010101";
		Trees_din <= x"ffda2691";
		wait for Clk_period;
		Addr <=  "00100101010110";
		Trees_din <= x"00612691";
		wait for Clk_period;
		Addr <=  "00100101010111";
		Trees_din <= x"0802c20c";
		wait for Clk_period;
		Addr <=  "00100101011000";
		Trees_din <= x"01146208";
		wait for Clk_period;
		Addr <=  "00100101011001";
		Trees_din <= x"0f03dc04";
		wait for Clk_period;
		Addr <=  "00100101011010";
		Trees_din <= x"00972691";
		wait for Clk_period;
		Addr <=  "00100101011011";
		Trees_din <= x"001d2691";
		wait for Clk_period;
		Addr <=  "00100101011100";
		Trees_din <= x"ffc32691";
		wait for Clk_period;
		Addr <=  "00100101011101";
		Trees_din <= x"1c002e04";
		wait for Clk_period;
		Addr <=  "00100101011110";
		Trees_din <= x"00622691";
		wait for Clk_period;
		Addr <=  "00100101011111";
		Trees_din <= x"0012b804";
		wait for Clk_period;
		Addr <=  "00100101100000";
		Trees_din <= x"ff762691";
		wait for Clk_period;
		Addr <=  "00100101100001";
		Trees_din <= x"fffc2691";
		wait for Clk_period;
		Addr <=  "00100101100010";
		Trees_din <= x"06f37f20";
		wait for Clk_period;
		Addr <=  "00100101100011";
		Trees_din <= x"04037810";
		wait for Clk_period;
		Addr <=  "00100101100100";
		Trees_din <= x"01107308";
		wait for Clk_period;
		Addr <=  "00100101100101";
		Trees_din <= x"13017904";
		wait for Clk_period;
		Addr <=  "00100101100110";
		Trees_din <= x"007a2691";
		wait for Clk_period;
		Addr <=  "00100101100111";
		Trees_din <= x"ffcb2691";
		wait for Clk_period;
		Addr <=  "00100101101000";
		Trees_din <= x"000d9f04";
		wait for Clk_period;
		Addr <=  "00100101101001";
		Trees_din <= x"ffab2691";
		wait for Clk_period;
		Addr <=  "00100101101010";
		Trees_din <= x"002a2691";
		wait for Clk_period;
		Addr <=  "00100101101011";
		Trees_din <= x"19009e08";
		wait for Clk_period;
		Addr <=  "00100101101100";
		Trees_din <= x"10055404";
		wait for Clk_period;
		Addr <=  "00100101101101";
		Trees_din <= x"ff812691";
		wait for Clk_period;
		Addr <=  "00100101101110";
		Trees_din <= x"fff32691";
		wait for Clk_period;
		Addr <=  "00100101101111";
		Trees_din <= x"0004c604";
		wait for Clk_period;
		Addr <=  "00100101110000";
		Trees_din <= x"ffd82691";
		wait for Clk_period;
		Addr <=  "00100101110001";
		Trees_din <= x"00632691";
		wait for Clk_period;
		Addr <=  "00100101110010";
		Trees_din <= x"001e7210";
		wait for Clk_period;
		Addr <=  "00100101110011";
		Trees_din <= x"09004808";
		wait for Clk_period;
		Addr <=  "00100101110100";
		Trees_din <= x"01081404";
		wait for Clk_period;
		Addr <=  "00100101110101";
		Trees_din <= x"00072691";
		wait for Clk_period;
		Addr <=  "00100101110110";
		Trees_din <= x"ff902691";
		wait for Clk_period;
		Addr <=  "00100101110111";
		Trees_din <= x"02062104";
		wait for Clk_period;
		Addr <=  "00100101111000";
		Trees_din <= x"fffe2691";
		wait for Clk_period;
		Addr <=  "00100101111001";
		Trees_din <= x"003f2691";
		wait for Clk_period;
		Addr <=  "00100101111010";
		Trees_din <= x"ff552691";
		wait for Clk_period;
		Addr <=  "00100101111011";
		Trees_din <= x"0207bf20";
		wait for Clk_period;
		Addr <=  "00100101111100";
		Trees_din <= x"06f5f210";
		wait for Clk_period;
		Addr <=  "00100101111101";
		Trees_din <= x"0900580c";
		wait for Clk_period;
		Addr <=  "00100101111110";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00100101111111";
		Trees_din <= x"00052691";
		wait for Clk_period;
		Addr <=  "00100110000000";
		Trees_din <= x"11028604";
		wait for Clk_period;
		Addr <=  "00100110000001";
		Trees_din <= x"ff432691";
		wait for Clk_period;
		Addr <=  "00100110000010";
		Trees_din <= x"ffe92691";
		wait for Clk_period;
		Addr <=  "00100110000011";
		Trees_din <= x"00352691";
		wait for Clk_period;
		Addr <=  "00100110000100";
		Trees_din <= x"0e01ce08";
		wait for Clk_period;
		Addr <=  "00100110000101";
		Trees_din <= x"1a00c604";
		wait for Clk_period;
		Addr <=  "00100110000110";
		Trees_din <= x"00812691";
		wait for Clk_period;
		Addr <=  "00100110000111";
		Trees_din <= x"fffa2691";
		wait for Clk_period;
		Addr <=  "00100110001000";
		Trees_din <= x"06f73b04";
		wait for Clk_period;
		Addr <=  "00100110001001";
		Trees_din <= x"fffd2691";
		wait for Clk_period;
		Addr <=  "00100110001010";
		Trees_din <= x"ff852691";
		wait for Clk_period;
		Addr <=  "00100110001011";
		Trees_din <= x"06f7891c";
		wait for Clk_period;
		Addr <=  "00100110001100";
		Trees_din <= x"04ff2e10";
		wait for Clk_period;
		Addr <=  "00100110001101";
		Trees_din <= x"02094408";
		wait for Clk_period;
		Addr <=  "00100110001110";
		Trees_din <= x"01117e04";
		wait for Clk_period;
		Addr <=  "00100110001111";
		Trees_din <= x"00722691";
		wait for Clk_period;
		Addr <=  "00100110010000";
		Trees_din <= x"ffe12691";
		wait for Clk_period;
		Addr <=  "00100110010001";
		Trees_din <= x"05f82b04";
		wait for Clk_period;
		Addr <=  "00100110010010";
		Trees_din <= x"00622691";
		wait for Clk_period;
		Addr <=  "00100110010011";
		Trees_din <= x"ffee2691";
		wait for Clk_period;
		Addr <=  "00100110010100";
		Trees_din <= x"0a034708";
		wait for Clk_period;
		Addr <=  "00100110010101";
		Trees_din <= x"00019004";
		wait for Clk_period;
		Addr <=  "00100110010110";
		Trees_din <= x"fffd2691";
		wait for Clk_period;
		Addr <=  "00100110010111";
		Trees_din <= x"ff702691";
		wait for Clk_period;
		Addr <=  "00100110011000";
		Trees_din <= x"00302691";
		wait for Clk_period;
		Addr <=  "00100110011001";
		Trees_din <= x"0afc8a10";
		wait for Clk_period;
		Addr <=  "00100110011010";
		Trees_din <= x"15009808";
		wait for Clk_period;
		Addr <=  "00100110011011";
		Trees_din <= x"0b041a04";
		wait for Clk_period;
		Addr <=  "00100110011100";
		Trees_din <= x"fff22691";
		wait for Clk_period;
		Addr <=  "00100110011101";
		Trees_din <= x"ffa32691";
		wait for Clk_period;
		Addr <=  "00100110011110";
		Trees_din <= x"1d004304";
		wait for Clk_period;
		Addr <=  "00100110011111";
		Trees_din <= x"001f2691";
		wait for Clk_period;
		Addr <=  "00100110100000";
		Trees_din <= x"00722691";
		wait for Clk_period;
		Addr <=  "00100110100001";
		Trees_din <= x"0802a504";
		wait for Clk_period;
		Addr <=  "00100110100010";
		Trees_din <= x"ff6a2691";
		wait for Clk_period;
		Addr <=  "00100110100011";
		Trees_din <= x"000e2691";
		wait for Clk_period;
		Addr <=  "00100110100100";
		Trees_din <= x"000b1e34";
		wait for Clk_period;
		Addr <=  "00100110100101";
		Trees_din <= x"03f85a08";
		wait for Clk_period;
		Addr <=  "00100110100110";
		Trees_din <= x"08031304";
		wait for Clk_period;
		Addr <=  "00100110100111";
		Trees_din <= x"ff82279d";
		wait for Clk_period;
		Addr <=  "00100110101000";
		Trees_din <= x"001c279d";
		wait for Clk_period;
		Addr <=  "00100110101001";
		Trees_din <= x"11fed318";
		wait for Clk_period;
		Addr <=  "00100110101010";
		Trees_din <= x"0e00d710";
		wait for Clk_period;
		Addr <=  "00100110101011";
		Trees_din <= x"0c035a08";
		wait for Clk_period;
		Addr <=  "00100110101100";
		Trees_din <= x"1f000004";
		wait for Clk_period;
		Addr <=  "00100110101101";
		Trees_din <= x"ff79279d";
		wait for Clk_period;
		Addr <=  "00100110101110";
		Trees_din <= x"001d279d";
		wait for Clk_period;
		Addr <=  "00100110101111";
		Trees_din <= x"17000004";
		wait for Clk_period;
		Addr <=  "00100110110000";
		Trees_din <= x"0068279d";
		wait for Clk_period;
		Addr <=  "00100110110001";
		Trees_din <= x"ffa6279d";
		wait for Clk_period;
		Addr <=  "00100110110010";
		Trees_din <= x"0c019a04";
		wait for Clk_period;
		Addr <=  "00100110110011";
		Trees_din <= x"005b279d";
		wait for Clk_period;
		Addr <=  "00100110110100";
		Trees_din <= x"0000279d";
		wait for Clk_period;
		Addr <=  "00100110110101";
		Trees_din <= x"0a046710";
		wait for Clk_period;
		Addr <=  "00100110110110";
		Trees_din <= x"13fdbb08";
		wait for Clk_period;
		Addr <=  "00100110110111";
		Trees_din <= x"0d00b304";
		wait for Clk_period;
		Addr <=  "00100110111000";
		Trees_din <= x"ffed279d";
		wait for Clk_period;
		Addr <=  "00100110111001";
		Trees_din <= x"0042279d";
		wait for Clk_period;
		Addr <=  "00100110111010";
		Trees_din <= x"0c004104";
		wait for Clk_period;
		Addr <=  "00100110111011";
		Trees_din <= x"0065279d";
		wait for Clk_period;
		Addr <=  "00100110111100";
		Trees_din <= x"ffe2279d";
		wait for Clk_period;
		Addr <=  "00100110111101";
		Trees_din <= x"0096279d";
		wait for Clk_period;
		Addr <=  "00100110111110";
		Trees_din <= x"18003620";
		wait for Clk_period;
		Addr <=  "00100110111111";
		Trees_din <= x"020db71c";
		wait for Clk_period;
		Addr <=  "00100111000000";
		Trees_din <= x"010db60c";
		wait for Clk_period;
		Addr <=  "00100111000001";
		Trees_din <= x"1d002d04";
		wait for Clk_period;
		Addr <=  "00100111000010";
		Trees_din <= x"fff3279d";
		wait for Clk_period;
		Addr <=  "00100111000011";
		Trees_din <= x"12fdea04";
		wait for Clk_period;
		Addr <=  "00100111000100";
		Trees_din <= x"000d279d";
		wait for Clk_period;
		Addr <=  "00100111000101";
		Trees_din <= x"00a2279d";
		wait for Clk_period;
		Addr <=  "00100111000110";
		Trees_din <= x"00115708";
		wait for Clk_period;
		Addr <=  "00100111000111";
		Trees_din <= x"0d00a704";
		wait for Clk_period;
		Addr <=  "00100111001000";
		Trees_din <= x"0045279d";
		wait for Clk_period;
		Addr <=  "00100111001001";
		Trees_din <= x"ff8f279d";
		wait for Clk_period;
		Addr <=  "00100111001010";
		Trees_din <= x"0c01b104";
		wait for Clk_period;
		Addr <=  "00100111001011";
		Trees_din <= x"0020279d";
		wait for Clk_period;
		Addr <=  "00100111001100";
		Trees_din <= x"0071279d";
		wait for Clk_period;
		Addr <=  "00100111001101";
		Trees_din <= x"ff9e279d";
		wait for Clk_period;
		Addr <=  "00100111001110";
		Trees_din <= x"1e005c14";
		wait for Clk_period;
		Addr <=  "00100111001111";
		Trees_din <= x"21000010";
		wait for Clk_period;
		Addr <=  "00100111010000";
		Trees_din <= x"08034308";
		wait for Clk_period;
		Addr <=  "00100111010001";
		Trees_din <= x"12fd8104";
		wait for Clk_period;
		Addr <=  "00100111010010";
		Trees_din <= x"006c279d";
		wait for Clk_period;
		Addr <=  "00100111010011";
		Trees_din <= x"ff9d279d";
		wait for Clk_period;
		Addr <=  "00100111010100";
		Trees_din <= x"1900ae04";
		wait for Clk_period;
		Addr <=  "00100111010101";
		Trees_din <= x"006d279d";
		wait for Clk_period;
		Addr <=  "00100111010110";
		Trees_din <= x"ffc7279d";
		wait for Clk_period;
		Addr <=  "00100111010111";
		Trees_din <= x"0089279d";
		wait for Clk_period;
		Addr <=  "00100111011000";
		Trees_din <= x"1a00d810";
		wait for Clk_period;
		Addr <=  "00100111011001";
		Trees_din <= x"10052908";
		wait for Clk_period;
		Addr <=  "00100111011010";
		Trees_din <= x"0afcd204";
		wait for Clk_period;
		Addr <=  "00100111011011";
		Trees_din <= x"ffdf279d";
		wait for Clk_period;
		Addr <=  "00100111011100";
		Trees_din <= x"000e279d";
		wait for Clk_period;
		Addr <=  "00100111011101";
		Trees_din <= x"03fe0704";
		wait for Clk_period;
		Addr <=  "00100111011110";
		Trees_din <= x"003a279d";
		wait for Clk_period;
		Addr <=  "00100111011111";
		Trees_din <= x"ff9a279d";
		wait for Clk_period;
		Addr <=  "00100111100000";
		Trees_din <= x"11fe7208";
		wait for Clk_period;
		Addr <=  "00100111100001";
		Trees_din <= x"1e005f04";
		wait for Clk_period;
		Addr <=  "00100111100010";
		Trees_din <= x"ff80279d";
		wait for Clk_period;
		Addr <=  "00100111100011";
		Trees_din <= x"fffe279d";
		wait for Clk_period;
		Addr <=  "00100111100100";
		Trees_din <= x"0e049504";
		wait for Clk_period;
		Addr <=  "00100111100101";
		Trees_din <= x"0068279d";
		wait for Clk_period;
		Addr <=  "00100111100110";
		Trees_din <= x"ffb3279d";
		wait for Clk_period;
		Addr <=  "00100111100111";
		Trees_din <= x"12028764";
		wait for Clk_period;
		Addr <=  "00100111101000";
		Trees_din <= x"06f37f34";
		wait for Clk_period;
		Addr <=  "00100111101001";
		Trees_din <= x"1200c318";
		wait for Clk_period;
		Addr <=  "00100111101010";
		Trees_din <= x"06f1460c";
		wait for Clk_period;
		Addr <=  "00100111101011";
		Trees_din <= x"000f9e04";
		wait for Clk_period;
		Addr <=  "00100111101100";
		Trees_din <= x"ff932909";
		wait for Clk_period;
		Addr <=  "00100111101101";
		Trees_din <= x"1a00b804";
		wait for Clk_period;
		Addr <=  "00100111101110";
		Trees_din <= x"ffc72909";
		wait for Clk_period;
		Addr <=  "00100111101111";
		Trees_din <= x"00522909";
		wait for Clk_period;
		Addr <=  "00100111110000";
		Trees_din <= x"1f000008";
		wait for Clk_period;
		Addr <=  "00100111110001";
		Trees_din <= x"0f03a804";
		wait for Clk_period;
		Addr <=  "00100111110010";
		Trees_din <= x"007a2909";
		wait for Clk_period;
		Addr <=  "00100111110011";
		Trees_din <= x"ffd42909";
		wait for Clk_period;
		Addr <=  "00100111110100";
		Trees_din <= x"ffa92909";
		wait for Clk_period;
		Addr <=  "00100111110101";
		Trees_din <= x"0207750c";
		wait for Clk_period;
		Addr <=  "00100111110110";
		Trees_din <= x"07005b08";
		wait for Clk_period;
		Addr <=  "00100111110111";
		Trees_din <= x"000d9f04";
		wait for Clk_period;
		Addr <=  "00100111111000";
		Trees_din <= x"fff32909";
		wait for Clk_period;
		Addr <=  "00100111111001";
		Trees_din <= x"007d2909";
		wait for Clk_period;
		Addr <=  "00100111111010";
		Trees_din <= x"ff912909";
		wait for Clk_period;
		Addr <=  "00100111111011";
		Trees_din <= x"0afaf208";
		wait for Clk_period;
		Addr <=  "00100111111100";
		Trees_din <= x"0f002c04";
		wait for Clk_period;
		Addr <=  "00100111111101";
		Trees_din <= x"00482909";
		wait for Clk_period;
		Addr <=  "00100111111110";
		Trees_din <= x"ffce2909";
		wait for Clk_period;
		Addr <=  "00100111111111";
		Trees_din <= x"05fdcb04";
		wait for Clk_period;
		Addr <=  "00101000000000";
		Trees_din <= x"ff7c2909";
		wait for Clk_period;
		Addr <=  "00101000000001";
		Trees_din <= x"00282909";
		wait for Clk_period;
		Addr <=  "00101000000010";
		Trees_din <= x"06f4631c";
		wait for Clk_period;
		Addr <=  "00101000000011";
		Trees_din <= x"12fdf60c";
		wait for Clk_period;
		Addr <=  "00101000000100";
		Trees_din <= x"0efe9604";
		wait for Clk_period;
		Addr <=  "00101000000101";
		Trees_din <= x"009b2909";
		wait for Clk_period;
		Addr <=  "00101000000110";
		Trees_din <= x"11fff404";
		wait for Clk_period;
		Addr <=  "00101000000111";
		Trees_din <= x"ff932909";
		wait for Clk_period;
		Addr <=  "00101000001000";
		Trees_din <= x"00322909";
		wait for Clk_period;
		Addr <=  "00101000001001";
		Trees_din <= x"010ad408";
		wait for Clk_period;
		Addr <=  "00101000001010";
		Trees_din <= x"11027704";
		wait for Clk_period;
		Addr <=  "00101000001011";
		Trees_din <= x"ffbd2909";
		wait for Clk_period;
		Addr <=  "00101000001100";
		Trees_din <= x"004d2909";
		wait for Clk_period;
		Addr <=  "00101000001101";
		Trees_din <= x"0012ed04";
		wait for Clk_period;
		Addr <=  "00101000001110";
		Trees_din <= x"ff6b2909";
		wait for Clk_period;
		Addr <=  "00101000001111";
		Trees_din <= x"fffa2909";
		wait for Clk_period;
		Addr <=  "00101000010000";
		Trees_din <= x"06f47704";
		wait for Clk_period;
		Addr <=  "00101000010001";
		Trees_din <= x"007b2909";
		wait for Clk_period;
		Addr <=  "00101000010010";
		Trees_din <= x"0d035b08";
		wait for Clk_period;
		Addr <=  "00101000010011";
		Trees_din <= x"09005b04";
		wait for Clk_period;
		Addr <=  "00101000010100";
		Trees_din <= x"fff92909";
		wait for Clk_period;
		Addr <=  "00101000010101";
		Trees_din <= x"ff9d2909";
		wait for Clk_period;
		Addr <=  "00101000010110";
		Trees_din <= x"0200e804";
		wait for Clk_period;
		Addr <=  "00101000010111";
		Trees_din <= x"ffc92909";
		wait for Clk_period;
		Addr <=  "00101000011000";
		Trees_din <= x"003c2909";
		wait for Clk_period;
		Addr <=  "00101000011001";
		Trees_din <= x"13013a20";
		wait for Clk_period;
		Addr <=  "00101000011010";
		Trees_din <= x"1c004214";
		wait for Clk_period;
		Addr <=  "00101000011011";
		Trees_din <= x"03033010";
		wait for Clk_period;
		Addr <=  "00101000011100";
		Trees_din <= x"0bf9c708";
		wait for Clk_period;
		Addr <=  "00101000011101";
		Trees_din <= x"0afb2604";
		wait for Clk_period;
		Addr <=  "00101000011110";
		Trees_din <= x"00552909";
		wait for Clk_period;
		Addr <=  "00101000011111";
		Trees_din <= x"ffc12909";
		wait for Clk_period;
		Addr <=  "00101000100000";
		Trees_din <= x"1c002b04";
		wait for Clk_period;
		Addr <=  "00101000100001";
		Trees_din <= x"00032909";
		wait for Clk_period;
		Addr <=  "00101000100010";
		Trees_din <= x"00812909";
		wait for Clk_period;
		Addr <=  "00101000100011";
		Trees_din <= x"ff8f2909";
		wait for Clk_period;
		Addr <=  "00101000100100";
		Trees_din <= x"1b004808";
		wait for Clk_period;
		Addr <=  "00101000100101";
		Trees_din <= x"0eff8004";
		wait for Clk_period;
		Addr <=  "00101000100110";
		Trees_din <= x"ff642909";
		wait for Clk_period;
		Addr <=  "00101000100111";
		Trees_din <= x"fffb2909";
		wait for Clk_period;
		Addr <=  "00101000101000";
		Trees_din <= x"00542909";
		wait for Clk_period;
		Addr <=  "00101000101001";
		Trees_din <= x"13016218";
		wait for Clk_period;
		Addr <=  "00101000101010";
		Trees_din <= x"06f50b08";
		wait for Clk_period;
		Addr <=  "00101000101011";
		Trees_din <= x"17005c04";
		wait for Clk_period;
		Addr <=  "00101000101100";
		Trees_din <= x"00652909";
		wait for Clk_period;
		Addr <=  "00101000101101";
		Trees_din <= x"ffe92909";
		wait for Clk_period;
		Addr <=  "00101000101110";
		Trees_din <= x"09005408";
		wait for Clk_period;
		Addr <=  "00101000101111";
		Trees_din <= x"0e040704";
		wait for Clk_period;
		Addr <=  "00101000110000";
		Trees_din <= x"ff8e2909";
		wait for Clk_period;
		Addr <=  "00101000110001";
		Trees_din <= x"005f2909";
		wait for Clk_period;
		Addr <=  "00101000110010";
		Trees_din <= x"01072b04";
		wait for Clk_period;
		Addr <=  "00101000110011";
		Trees_din <= x"ffd12909";
		wait for Clk_period;
		Addr <=  "00101000110100";
		Trees_din <= x"ff332909";
		wait for Clk_period;
		Addr <=  "00101000110101";
		Trees_din <= x"00111710";
		wait for Clk_period;
		Addr <=  "00101000110110";
		Trees_din <= x"1b003808";
		wait for Clk_period;
		Addr <=  "00101000110111";
		Trees_din <= x"1f000004";
		wait for Clk_period;
		Addr <=  "00101000111000";
		Trees_din <= x"ff8d2909";
		wait for Clk_period;
		Addr <=  "00101000111001";
		Trees_din <= x"002d2909";
		wait for Clk_period;
		Addr <=  "00101000111010";
		Trees_din <= x"18004904";
		wait for Clk_period;
		Addr <=  "00101000111011";
		Trees_din <= x"00502909";
		wait for Clk_period;
		Addr <=  "00101000111100";
		Trees_din <= x"ffd12909";
		wait for Clk_period;
		Addr <=  "00101000111101";
		Trees_din <= x"08005c08";
		wait for Clk_period;
		Addr <=  "00101000111110";
		Trees_din <= x"11043804";
		wait for Clk_period;
		Addr <=  "00101000111111";
		Trees_din <= x"00712909";
		wait for Clk_period;
		Addr <=  "00101001000000";
		Trees_din <= x"ff842909";
		wait for Clk_period;
		Addr <=  "00101001000001";
		Trees_din <= x"00932909";
		wait for Clk_period;
		Addr <=  "00101001000010";
		Trees_din <= x"09005e74";
		wait for Clk_period;
		Addr <=  "00101001000011";
		Trees_din <= x"05fc2238";
		wait for Clk_period;
		Addr <=  "00101001000100";
		Trees_din <= x"1d004418";
		wait for Clk_period;
		Addr <=  "00101001000101";
		Trees_din <= x"05fc0a10";
		wait for Clk_period;
		Addr <=  "00101001000110";
		Trees_din <= x"1a00de08";
		wait for Clk_period;
		Addr <=  "00101001000111";
		Trees_din <= x"0afaca04";
		wait for Clk_period;
		Addr <=  "00101001001000";
		Trees_din <= x"ffc829fd";
		wait for Clk_period;
		Addr <=  "00101001001001";
		Trees_din <= x"003929fd";
		wait for Clk_period;
		Addr <=  "00101001001010";
		Trees_din <= x"0f00a304";
		wait for Clk_period;
		Addr <=  "00101001001011";
		Trees_din <= x"ffce29fd";
		wait for Clk_period;
		Addr <=  "00101001001100";
		Trees_din <= x"001329fd";
		wait for Clk_period;
		Addr <=  "00101001001101";
		Trees_din <= x"07005304";
		wait for Clk_period;
		Addr <=  "00101001001110";
		Trees_din <= x"001729fd";
		wait for Clk_period;
		Addr <=  "00101001001111";
		Trees_din <= x"ff4429fd";
		wait for Clk_period;
		Addr <=  "00101001010000";
		Trees_din <= x"06f56510";
		wait for Clk_period;
		Addr <=  "00101001010001";
		Trees_din <= x"06f33608";
		wait for Clk_period;
		Addr <=  "00101001010010";
		Trees_din <= x"04037804";
		wait for Clk_period;
		Addr <=  "00101001010011";
		Trees_din <= x"000f29fd";
		wait for Clk_period;
		Addr <=  "00101001010100";
		Trees_din <= x"ff8729fd";
		wait for Clk_period;
		Addr <=  "00101001010101";
		Trees_din <= x"15008904";
		wait for Clk_period;
		Addr <=  "00101001010110";
		Trees_din <= x"000029fd";
		wait for Clk_period;
		Addr <=  "00101001010111";
		Trees_din <= x"ff9129fd";
		wait for Clk_period;
		Addr <=  "00101001011000";
		Trees_din <= x"0c01f408";
		wait for Clk_period;
		Addr <=  "00101001011001";
		Trees_din <= x"1d004904";
		wait for Clk_period;
		Addr <=  "00101001011010";
		Trees_din <= x"ffa229fd";
		wait for Clk_period;
		Addr <=  "00101001011011";
		Trees_din <= x"000729fd";
		wait for Clk_period;
		Addr <=  "00101001011100";
		Trees_din <= x"010e0804";
		wait for Clk_period;
		Addr <=  "00101001011101";
		Trees_din <= x"000229fd";
		wait for Clk_period;
		Addr <=  "00101001011110";
		Trees_din <= x"007329fd";
		wait for Clk_period;
		Addr <=  "00101001011111";
		Trees_din <= x"06f54920";
		wait for Clk_period;
		Addr <=  "00101001100000";
		Trees_din <= x"06f45810";
		wait for Clk_period;
		Addr <=  "00101001100001";
		Trees_din <= x"06f36508";
		wait for Clk_period;
		Addr <=  "00101001100010";
		Trees_din <= x"0c01b504";
		wait for Clk_period;
		Addr <=  "00101001100011";
		Trees_din <= x"ffe929fd";
		wait for Clk_period;
		Addr <=  "00101001100100";
		Trees_din <= x"006929fd";
		wait for Clk_period;
		Addr <=  "00101001100101";
		Trees_din <= x"12015404";
		wait for Clk_period;
		Addr <=  "00101001100110";
		Trees_din <= x"ff8929fd";
		wait for Clk_period;
		Addr <=  "00101001100111";
		Trees_din <= x"000a29fd";
		wait for Clk_period;
		Addr <=  "00101001101000";
		Trees_din <= x"10052108";
		wait for Clk_period;
		Addr <=  "00101001101001";
		Trees_din <= x"0100f904";
		wait for Clk_period;
		Addr <=  "00101001101010";
		Trees_din <= x"000029fd";
		wait for Clk_period;
		Addr <=  "00101001101011";
		Trees_din <= x"00a829fd";
		wait for Clk_period;
		Addr <=  "00101001101100";
		Trees_din <= x"13ffc104";
		wait for Clk_period;
		Addr <=  "00101001101101";
		Trees_din <= x"ffae29fd";
		wait for Clk_period;
		Addr <=  "00101001101110";
		Trees_din <= x"004c29fd";
		wait for Clk_period;
		Addr <=  "00101001101111";
		Trees_din <= x"0afac20c";
		wait for Clk_period;
		Addr <=  "00101001110000";
		Trees_din <= x"05ffdf08";
		wait for Clk_period;
		Addr <=  "00101001110001";
		Trees_din <= x"00087804";
		wait for Clk_period;
		Addr <=  "00101001110010";
		Trees_din <= x"000829fd";
		wait for Clk_period;
		Addr <=  "00101001110011";
		Trees_din <= x"009c29fd";
		wait for Clk_period;
		Addr <=  "00101001110100";
		Trees_din <= x"ffa729fd";
		wait for Clk_period;
		Addr <=  "00101001110101";
		Trees_din <= x"1d004508";
		wait for Clk_period;
		Addr <=  "00101001110110";
		Trees_din <= x"08033204";
		wait for Clk_period;
		Addr <=  "00101001110111";
		Trees_din <= x"ffc129fd";
		wait for Clk_period;
		Addr <=  "00101001111000";
		Trees_din <= x"004029fd";
		wait for Clk_period;
		Addr <=  "00101001111001";
		Trees_din <= x"18004604";
		wait for Clk_period;
		Addr <=  "00101001111010";
		Trees_din <= x"004e29fd";
		wait for Clk_period;
		Addr <=  "00101001111011";
		Trees_din <= x"ffef29fd";
		wait for Clk_period;
		Addr <=  "00101001111100";
		Trees_din <= x"0f002404";
		wait for Clk_period;
		Addr <=  "00101001111101";
		Trees_din <= x"000e29fd";
		wait for Clk_period;
		Addr <=  "00101001111110";
		Trees_din <= x"007029fd";
		wait for Clk_period;
		Addr <=  "00101001111111";
		Trees_din <= x"09005e70";
		wait for Clk_period;
		Addr <=  "00101010000000";
		Trees_din <= x"000f6f3c";
		wait for Clk_period;
		Addr <=  "00101010000001";
		Trees_din <= x"0c014020";
		wait for Clk_period;
		Addr <=  "00101010000010";
		Trees_din <= x"06f65a10";
		wait for Clk_period;
		Addr <=  "00101010000011";
		Trees_din <= x"0af7c608";
		wait for Clk_period;
		Addr <=  "00101010000100";
		Trees_din <= x"13fda304";
		wait for Clk_period;
		Addr <=  "00101010000101";
		Trees_din <= x"000a2ae9";
		wait for Clk_period;
		Addr <=  "00101010000110";
		Trees_din <= x"ff6a2ae9";
		wait for Clk_period;
		Addr <=  "00101010000111";
		Trees_din <= x"05fe4a04";
		wait for Clk_period;
		Addr <=  "00101010001000";
		Trees_din <= x"001c2ae9";
		wait for Clk_period;
		Addr <=  "00101010001001";
		Trees_din <= x"ff7b2ae9";
		wait for Clk_period;
		Addr <=  "00101010001010";
		Trees_din <= x"01029908";
		wait for Clk_period;
		Addr <=  "00101010001011";
		Trees_din <= x"05ff3504";
		wait for Clk_period;
		Addr <=  "00101010001100";
		Trees_din <= x"002b2ae9";
		wait for Clk_period;
		Addr <=  "00101010001101";
		Trees_din <= x"ff9c2ae9";
		wait for Clk_period;
		Addr <=  "00101010001110";
		Trees_din <= x"0e045004";
		wait for Clk_period;
		Addr <=  "00101010001111";
		Trees_din <= x"ff8e2ae9";
		wait for Clk_period;
		Addr <=  "00101010010000";
		Trees_din <= x"003e2ae9";
		wait for Clk_period;
		Addr <=  "00101010010001";
		Trees_din <= x"05f88b0c";
		wait for Clk_period;
		Addr <=  "00101010010010";
		Trees_din <= x"0ef9a904";
		wait for Clk_period;
		Addr <=  "00101010010011";
		Trees_din <= x"00472ae9";
		wait for Clk_period;
		Addr <=  "00101010010100";
		Trees_din <= x"1a00f904";
		wait for Clk_period;
		Addr <=  "00101010010101";
		Trees_din <= x"ff7b2ae9";
		wait for Clk_period;
		Addr <=  "00101010010110";
		Trees_din <= x"00002ae9";
		wait for Clk_period;
		Addr <=  "00101010010111";
		Trees_din <= x"05f8d108";
		wait for Clk_period;
		Addr <=  "00101010011000";
		Trees_din <= x"09005104";
		wait for Clk_period;
		Addr <=  "00101010011001";
		Trees_din <= x"00d42ae9";
		wait for Clk_period;
		Addr <=  "00101010011010";
		Trees_din <= x"00112ae9";
		wait for Clk_period;
		Addr <=  "00101010011011";
		Trees_din <= x"010a1f04";
		wait for Clk_period;
		Addr <=  "00101010011100";
		Trees_din <= x"00162ae9";
		wait for Clk_period;
		Addr <=  "00101010011101";
		Trees_din <= x"ffe32ae9";
		wait for Clk_period;
		Addr <=  "00101010011110";
		Trees_din <= x"1603a620";
		wait for Clk_period;
		Addr <=  "00101010011111";
		Trees_din <= x"18003b10";
		wait for Clk_period;
		Addr <=  "00101010100000";
		Trees_din <= x"0f016808";
		wait for Clk_period;
		Addr <=  "00101010100001";
		Trees_din <= x"1700f604";
		wait for Clk_period;
		Addr <=  "00101010100010";
		Trees_din <= x"00492ae9";
		wait for Clk_period;
		Addr <=  "00101010100011";
		Trees_din <= x"ffae2ae9";
		wait for Clk_period;
		Addr <=  "00101010100100";
		Trees_din <= x"1f000c04";
		wait for Clk_period;
		Addr <=  "00101010100101";
		Trees_din <= x"008d2ae9";
		wait for Clk_period;
		Addr <=  "00101010100110";
		Trees_din <= x"ffd32ae9";
		wait for Clk_period;
		Addr <=  "00101010100111";
		Trees_din <= x"1b003608";
		wait for Clk_period;
		Addr <=  "00101010101000";
		Trees_din <= x"06f4ad04";
		wait for Clk_period;
		Addr <=  "00101010101001";
		Trees_din <= x"00562ae9";
		wait for Clk_period;
		Addr <=  "00101010101010";
		Trees_din <= x"ff982ae9";
		wait for Clk_period;
		Addr <=  "00101010101011";
		Trees_din <= x"02071404";
		wait for Clk_period;
		Addr <=  "00101010101100";
		Trees_din <= x"00272ae9";
		wait for Clk_period;
		Addr <=  "00101010101101";
		Trees_din <= x"ffd42ae9";
		wait for Clk_period;
		Addr <=  "00101010101110";
		Trees_din <= x"03f7e310";
		wait for Clk_period;
		Addr <=  "00101010101111";
		Trees_din <= x"0f000708";
		wait for Clk_period;
		Addr <=  "00101010110000";
		Trees_din <= x"19008904";
		wait for Clk_period;
		Addr <=  "00101010110001";
		Trees_din <= x"005b2ae9";
		wait for Clk_period;
		Addr <=  "00101010110010";
		Trees_din <= x"ffa02ae9";
		wait for Clk_period;
		Addr <=  "00101010110011";
		Trees_din <= x"04f9a004";
		wait for Clk_period;
		Addr <=  "00101010110100";
		Trees_din <= x"00522ae9";
		wait for Clk_period;
		Addr <=  "00101010110101";
		Trees_din <= x"ffdf2ae9";
		wait for Clk_period;
		Addr <=  "00101010110110";
		Trees_din <= x"00952ae9";
		wait for Clk_period;
		Addr <=  "00101010110111";
		Trees_din <= x"010a4204";
		wait for Clk_period;
		Addr <=  "00101010111000";
		Trees_din <= x"001a2ae9";
		wait for Clk_period;
		Addr <=  "00101010111001";
		Trees_din <= x"00732ae9";
		wait for Clk_period;
		Addr <=  "00101010111010";
		Trees_din <= x"0003aa34";
		wait for Clk_period;
		Addr <=  "00101010111011";
		Trees_din <= x"1b003d18";
		wait for Clk_period;
		Addr <=  "00101010111100";
		Trees_din <= x"1f000010";
		wait for Clk_period;
		Addr <=  "00101010111101";
		Trees_din <= x"08023808";
		wait for Clk_period;
		Addr <=  "00101010111110";
		Trees_din <= x"10f99904";
		wait for Clk_period;
		Addr <=  "00101010111111";
		Trees_din <= x"ffd92c35";
		wait for Clk_period;
		Addr <=  "00101011000000";
		Trees_din <= x"ff7b2c35";
		wait for Clk_period;
		Addr <=  "00101011000001";
		Trees_din <= x"08029604";
		wait for Clk_period;
		Addr <=  "00101011000010";
		Trees_din <= x"00492c35";
		wait for Clk_period;
		Addr <=  "00101011000011";
		Trees_din <= x"ffa02c35";
		wait for Clk_period;
		Addr <=  "00101011000100";
		Trees_din <= x"07005304";
		wait for Clk_period;
		Addr <=  "00101011000101";
		Trees_din <= x"00442c35";
		wait for Clk_period;
		Addr <=  "00101011000110";
		Trees_din <= x"ffcb2c35";
		wait for Clk_period;
		Addr <=  "00101011000111";
		Trees_din <= x"07005814";
		wait for Clk_period;
		Addr <=  "00101011001000";
		Trees_din <= x"0c01fd0c";
		wait for Clk_period;
		Addr <=  "00101011001001";
		Trees_din <= x"0c012008";
		wait for Clk_period;
		Addr <=  "00101011001010";
		Trees_din <= x"13fdce04";
		wait for Clk_period;
		Addr <=  "00101011001011";
		Trees_din <= x"001b2c35";
		wait for Clk_period;
		Addr <=  "00101011001100";
		Trees_din <= x"ffcf2c35";
		wait for Clk_period;
		Addr <=  "00101011001101";
		Trees_din <= x"007d2c35";
		wait for Clk_period;
		Addr <=  "00101011001110";
		Trees_din <= x"1102d204";
		wait for Clk_period;
		Addr <=  "00101011001111";
		Trees_din <= x"ffa72c35";
		wait for Clk_period;
		Addr <=  "00101011010000";
		Trees_din <= x"00272c35";
		wait for Clk_period;
		Addr <=  "00101011010001";
		Trees_din <= x"1c003504";
		wait for Clk_period;
		Addr <=  "00101011010010";
		Trees_din <= x"00122c35";
		wait for Clk_period;
		Addr <=  "00101011010011";
		Trees_din <= x"ff972c35";
		wait for Clk_period;
		Addr <=  "00101011010100";
		Trees_din <= x"02ffbf34";
		wait for Clk_period;
		Addr <=  "00101011010101";
		Trees_din <= x"06f68b14";
		wait for Clk_period;
		Addr <=  "00101011010110";
		Trees_din <= x"0bf95304";
		wait for Clk_period;
		Addr <=  "00101011010111";
		Trees_din <= x"ffbf2c35";
		wait for Clk_period;
		Addr <=  "00101011011000";
		Trees_din <= x"1c003e08";
		wait for Clk_period;
		Addr <=  "00101011011001";
		Trees_din <= x"10f95704";
		wait for Clk_period;
		Addr <=  "00101011011010";
		Trees_din <= x"00042c35";
		wait for Clk_period;
		Addr <=  "00101011011011";
		Trees_din <= x"008b2c35";
		wait for Clk_period;
		Addr <=  "00101011011100";
		Trees_din <= x"13fe2d04";
		wait for Clk_period;
		Addr <=  "00101011011101";
		Trees_din <= x"ffae2c35";
		wait for Clk_period;
		Addr <=  "00101011011110";
		Trees_din <= x"00452c35";
		wait for Clk_period;
		Addr <=  "00101011011111";
		Trees_din <= x"0f003e10";
		wait for Clk_period;
		Addr <=  "00101011100000";
		Trees_din <= x"00090508";
		wait for Clk_period;
		Addr <=  "00101011100001";
		Trees_din <= x"01012e04";
		wait for Clk_period;
		Addr <=  "00101011100010";
		Trees_din <= x"00352c35";
		wait for Clk_period;
		Addr <=  "00101011100011";
		Trees_din <= x"ffb92c35";
		wait for Clk_period;
		Addr <=  "00101011100100";
		Trees_din <= x"0a02bd04";
		wait for Clk_period;
		Addr <=  "00101011100101";
		Trees_din <= x"00862c35";
		wait for Clk_period;
		Addr <=  "00101011100110";
		Trees_din <= x"00142c35";
		wait for Clk_period;
		Addr <=  "00101011100111";
		Trees_din <= x"07005a08";
		wait for Clk_period;
		Addr <=  "00101011101000";
		Trees_din <= x"07005804";
		wait for Clk_period;
		Addr <=  "00101011101001";
		Trees_din <= x"00112c35";
		wait for Clk_period;
		Addr <=  "00101011101010";
		Trees_din <= x"ff882c35";
		wait for Clk_period;
		Addr <=  "00101011101011";
		Trees_din <= x"0afd0d04";
		wait for Clk_period;
		Addr <=  "00101011101100";
		Trees_din <= x"00012c35";
		wait for Clk_period;
		Addr <=  "00101011101101";
		Trees_din <= x"005f2c35";
		wait for Clk_period;
		Addr <=  "00101011101110";
		Trees_din <= x"0200c420";
		wait for Clk_period;
		Addr <=  "00101011101111";
		Trees_din <= x"06f6f110";
		wait for Clk_period;
		Addr <=  "00101011110000";
		Trees_din <= x"20040008";
		wait for Clk_period;
		Addr <=  "00101011110001";
		Trees_din <= x"1d004f04";
		wait for Clk_period;
		Addr <=  "00101011110010";
		Trees_din <= x"00512c35";
		wait for Clk_period;
		Addr <=  "00101011110011";
		Trees_din <= x"ffa52c35";
		wait for Clk_period;
		Addr <=  "00101011110100";
		Trees_din <= x"1701d504";
		wait for Clk_period;
		Addr <=  "00101011110101";
		Trees_din <= x"ff5d2c35";
		wait for Clk_period;
		Addr <=  "00101011110110";
		Trees_din <= x"ffef2c35";
		wait for Clk_period;
		Addr <=  "00101011110111";
		Trees_din <= x"10047f08";
		wait for Clk_period;
		Addr <=  "00101011111000";
		Trees_din <= x"00090504";
		wait for Clk_period;
		Addr <=  "00101011111001";
		Trees_din <= x"ffcd2c35";
		wait for Clk_period;
		Addr <=  "00101011111010";
		Trees_din <= x"008b2c35";
		wait for Clk_period;
		Addr <=  "00101011111011";
		Trees_din <= x"01050204";
		wait for Clk_period;
		Addr <=  "00101011111100";
		Trees_din <= x"00412c35";
		wait for Clk_period;
		Addr <=  "00101011111101";
		Trees_din <= x"ff882c35";
		wait for Clk_period;
		Addr <=  "00101011111110";
		Trees_din <= x"0d037b10";
		wait for Clk_period;
		Addr <=  "00101011111111";
		Trees_din <= x"1402f408";
		wait for Clk_period;
		Addr <=  "00101100000000";
		Trees_din <= x"1603ae04";
		wait for Clk_period;
		Addr <=  "00101100000001";
		Trees_din <= x"ffe22c35";
		wait for Clk_period;
		Addr <=  "00101100000010";
		Trees_din <= x"00122c35";
		wait for Clk_period;
		Addr <=  "00101100000011";
		Trees_din <= x"1403b404";
		wait for Clk_period;
		Addr <=  "00101100000100";
		Trees_din <= x"00412c35";
		wait for Clk_period;
		Addr <=  "00101100000101";
		Trees_din <= x"fff22c35";
		wait for Clk_period;
		Addr <=  "00101100000110";
		Trees_din <= x"02072e08";
		wait for Clk_period;
		Addr <=  "00101100000111";
		Trees_din <= x"1700de04";
		wait for Clk_period;
		Addr <=  "00101100001000";
		Trees_din <= x"00502c35";
		wait for Clk_period;
		Addr <=  "00101100001001";
		Trees_din <= x"fff22c35";
		wait for Clk_period;
		Addr <=  "00101100001010";
		Trees_din <= x"03f94d04";
		wait for Clk_period;
		Addr <=  "00101100001011";
		Trees_din <= x"001e2c35";
		wait for Clk_period;
		Addr <=  "00101100001100";
		Trees_din <= x"ff702c35";
		wait for Clk_period;
		Addr <=  "00101100001101";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00101100001110";
		Trees_din <= x"09005e64";
		wait for Clk_period;
		Addr <=  "00101100001111";
		Trees_din <= x"05fc2224";
		wait for Clk_period;
		Addr <=  "00101100010000";
		Trees_din <= x"10f71004";
		wait for Clk_period;
		Addr <=  "00101100010001";
		Trees_din <= x"006c2d0d";
		wait for Clk_period;
		Addr <=  "00101100010010";
		Trees_din <= x"0af7c610";
		wait for Clk_period;
		Addr <=  "00101100010011";
		Trees_din <= x"03f79308";
		wait for Clk_period;
		Addr <=  "00101100010100";
		Trees_din <= x"0203b004";
		wait for Clk_period;
		Addr <=  "00101100010101";
		Trees_din <= x"ffd12d0d";
		wait for Clk_period;
		Addr <=  "00101100010110";
		Trees_din <= x"00652d0d";
		wait for Clk_period;
		Addr <=  "00101100010111";
		Trees_din <= x"0b03e304";
		wait for Clk_period;
		Addr <=  "00101100011000";
		Trees_din <= x"00132d0d";
		wait for Clk_period;
		Addr <=  "00101100011001";
		Trees_din <= x"ff752d0d";
		wait for Clk_period;
		Addr <=  "00101100011010";
		Trees_din <= x"0af7e808";
		wait for Clk_period;
		Addr <=  "00101100011011";
		Trees_din <= x"1703d804";
		wait for Clk_period;
		Addr <=  "00101100011100";
		Trees_din <= x"007e2d0d";
		wait for Clk_period;
		Addr <=  "00101100011101";
		Trees_din <= x"ffe12d0d";
		wait for Clk_period;
		Addr <=  "00101100011110";
		Trees_din <= x"0afaca04";
		wait for Clk_period;
		Addr <=  "00101100011111";
		Trees_din <= x"ffb92d0d";
		wait for Clk_period;
		Addr <=  "00101100100000";
		Trees_din <= x"fffd2d0d";
		wait for Clk_period;
		Addr <=  "00101100100001";
		Trees_din <= x"06f54920";
		wait for Clk_period;
		Addr <=  "00101100100010";
		Trees_din <= x"06f45810";
		wait for Clk_period;
		Addr <=  "00101100100011";
		Trees_din <= x"000f6f08";
		wait for Clk_period;
		Addr <=  "00101100100100";
		Trees_din <= x"05fc4404";
		wait for Clk_period;
		Addr <=  "00101100100101";
		Trees_din <= x"005a2d0d";
		wait for Clk_period;
		Addr <=  "00101100100110";
		Trees_din <= x"ffbf2d0d";
		wait for Clk_period;
		Addr <=  "00101100100111";
		Trees_din <= x"16035e04";
		wait for Clk_period;
		Addr <=  "00101100101000";
		Trees_din <= x"00732d0d";
		wait for Clk_period;
		Addr <=  "00101100101001";
		Trees_din <= x"ffec2d0d";
		wait for Clk_period;
		Addr <=  "00101100101010";
		Trees_din <= x"020abe08";
		wait for Clk_period;
		Addr <=  "00101100101011";
		Trees_din <= x"11fe1b04";
		wait for Clk_period;
		Addr <=  "00101100101100";
		Trees_din <= x"ffec2d0d";
		wait for Clk_period;
		Addr <=  "00101100101101";
		Trees_din <= x"00942d0d";
		wait for Clk_period;
		Addr <=  "00101100101110";
		Trees_din <= x"09005804";
		wait for Clk_period;
		Addr <=  "00101100101111";
		Trees_din <= x"ffb42d0d";
		wait for Clk_period;
		Addr <=  "00101100110000";
		Trees_din <= x"00482d0d";
		wait for Clk_period;
		Addr <=  "00101100110001";
		Trees_din <= x"0a01b510";
		wait for Clk_period;
		Addr <=  "00101100110010";
		Trees_din <= x"1b003b08";
		wait for Clk_period;
		Addr <=  "00101100110011";
		Trees_din <= x"0102bb04";
		wait for Clk_period;
		Addr <=  "00101100110100";
		Trees_din <= x"00202d0d";
		wait for Clk_period;
		Addr <=  "00101100110101";
		Trees_din <= x"ffcd2d0d";
		wait for Clk_period;
		Addr <=  "00101100110110";
		Trees_din <= x"0500cb04";
		wait for Clk_period;
		Addr <=  "00101100110111";
		Trees_din <= x"004b2d0d";
		wait for Clk_period;
		Addr <=  "00101100111000";
		Trees_din <= x"ffbb2d0d";
		wait for Clk_period;
		Addr <=  "00101100111001";
		Trees_din <= x"08032b08";
		wait for Clk_period;
		Addr <=  "00101100111010";
		Trees_din <= x"000f6f04";
		wait for Clk_period;
		Addr <=  "00101100111011";
		Trees_din <= x"ffa52d0d";
		wait for Clk_period;
		Addr <=  "00101100111100";
		Trees_din <= x"00032d0d";
		wait for Clk_period;
		Addr <=  "00101100111101";
		Trees_din <= x"09005704";
		wait for Clk_period;
		Addr <=  "00101100111110";
		Trees_din <= x"00672d0d";
		wait for Clk_period;
		Addr <=  "00101100111111";
		Trees_din <= x"ffbc2d0d";
		wait for Clk_period;
		Addr <=  "00101101000000";
		Trees_din <= x"010a4204";
		wait for Clk_period;
		Addr <=  "00101101000001";
		Trees_din <= x"001a2d0d";
		wait for Clk_period;
		Addr <=  "00101101000010";
		Trees_din <= x"006f2d0d";
		wait for Clk_period;
		Addr <=  "00101101000011";
		Trees_din <= x"0003aa2c";
		wait for Clk_period;
		Addr <=  "00101101000100";
		Trees_din <= x"09005418";
		wait for Clk_period;
		Addr <=  "00101101000101";
		Trees_din <= x"1e006108";
		wait for Clk_period;
		Addr <=  "00101101000110";
		Trees_din <= x"1c002404";
		wait for Clk_period;
		Addr <=  "00101101000111";
		Trees_din <= x"00142db1";
		wait for Clk_period;
		Addr <=  "00101101001000";
		Trees_din <= x"ff912db1";
		wait for Clk_period;
		Addr <=  "00101101001001";
		Trees_din <= x"1004380c";
		wait for Clk_period;
		Addr <=  "00101101001010";
		Trees_din <= x"19008604";
		wait for Clk_period;
		Addr <=  "00101101001011";
		Trees_din <= x"ffcf2db1";
		wait for Clk_period;
		Addr <=  "00101101001100";
		Trees_din <= x"0bff0b04";
		wait for Clk_period;
		Addr <=  "00101101001101";
		Trees_din <= x"00192db1";
		wait for Clk_period;
		Addr <=  "00101101001110";
		Trees_din <= x"007a2db1";
		wait for Clk_period;
		Addr <=  "00101101001111";
		Trees_din <= x"ffab2db1";
		wait for Clk_period;
		Addr <=  "00101101010000";
		Trees_din <= x"15008708";
		wait for Clk_period;
		Addr <=  "00101101010001";
		Trees_din <= x"05fd3d04";
		wait for Clk_period;
		Addr <=  "00101101010010";
		Trees_din <= x"ffe42db1";
		wait for Clk_period;
		Addr <=  "00101101010011";
		Trees_din <= x"00572db1";
		wait for Clk_period;
		Addr <=  "00101101010100";
		Trees_din <= x"15009b04";
		wait for Clk_period;
		Addr <=  "00101101010101";
		Trees_din <= x"ff7c2db1";
		wait for Clk_period;
		Addr <=  "00101101010110";
		Trees_din <= x"14023404";
		wait for Clk_period;
		Addr <=  "00101101010111";
		Trees_din <= x"ffaa2db1";
		wait for Clk_period;
		Addr <=  "00101101011000";
		Trees_din <= x"00222db1";
		wait for Clk_period;
		Addr <=  "00101101011001";
		Trees_din <= x"02fdcd10";
		wait for Clk_period;
		Addr <=  "00101101011010";
		Trees_din <= x"0108bd08";
		wait for Clk_period;
		Addr <=  "00101101011011";
		Trees_din <= x"00054504";
		wait for Clk_period;
		Addr <=  "00101101011100";
		Trees_din <= x"00052db1";
		wait for Clk_period;
		Addr <=  "00101101011101";
		Trees_din <= x"00782db1";
		wait for Clk_period;
		Addr <=  "00101101011110";
		Trees_din <= x"0f00ba04";
		wait for Clk_period;
		Addr <=  "00101101011111";
		Trees_din <= x"00302db1";
		wait for Clk_period;
		Addr <=  "00101101100000";
		Trees_din <= x"ffc22db1";
		wait for Clk_period;
		Addr <=  "00101101100001";
		Trees_din <= x"0306c214";
		wait for Clk_period;
		Addr <=  "00101101100010";
		Trees_din <= x"09005e10";
		wait for Clk_period;
		Addr <=  "00101101100011";
		Trees_din <= x"18004808";
		wait for Clk_period;
		Addr <=  "00101101100100";
		Trees_din <= x"1b003804";
		wait for Clk_period;
		Addr <=  "00101101100101";
		Trees_din <= x"fffb2db1";
		wait for Clk_period;
		Addr <=  "00101101100110";
		Trees_din <= x"00192db1";
		wait for Clk_period;
		Addr <=  "00101101100111";
		Trees_din <= x"1b003f04";
		wait for Clk_period;
		Addr <=  "00101101101000";
		Trees_din <= x"ffac2db1";
		wait for Clk_period;
		Addr <=  "00101101101001";
		Trees_din <= x"00032db1";
		wait for Clk_period;
		Addr <=  "00101101101010";
		Trees_din <= x"005d2db1";
		wait for Clk_period;
		Addr <=  "00101101101011";
		Trees_din <= x"ff982db1";
		wait for Clk_period;
		Addr <=  "00101101101100";
		Trees_din <= x"0003aa28";
		wait for Clk_period;
		Addr <=  "00101101101101";
		Trees_din <= x"11010008";
		wait for Clk_period;
		Addr <=  "00101101101110";
		Trees_din <= x"0f03a304";
		wait for Clk_period;
		Addr <=  "00101101101111";
		Trees_din <= x"ff872ead";
		wait for Clk_period;
		Addr <=  "00101101110000";
		Trees_din <= x"000c2ead";
		wait for Clk_period;
		Addr <=  "00101101110001";
		Trees_din <= x"02006c0c";
		wait for Clk_period;
		Addr <=  "00101101110010";
		Trees_din <= x"02fba504";
		wait for Clk_period;
		Addr <=  "00101101110011";
		Trees_din <= x"00272ead";
		wait for Clk_period;
		Addr <=  "00101101110100";
		Trees_din <= x"0bf96b04";
		wait for Clk_period;
		Addr <=  "00101101110101";
		Trees_din <= x"fff12ead";
		wait for Clk_period;
		Addr <=  "00101101110110";
		Trees_din <= x"ff872ead";
		wait for Clk_period;
		Addr <=  "00101101110111";
		Trees_din <= x"0204540c";
		wait for Clk_period;
		Addr <=  "00101101111000";
		Trees_din <= x"05fd9808";
		wait for Clk_period;
		Addr <=  "00101101111001";
		Trees_din <= x"09005604";
		wait for Clk_period;
		Addr <=  "00101101111010";
		Trees_din <= x"00772ead";
		wait for Clk_period;
		Addr <=  "00101101111011";
		Trees_din <= x"ffeb2ead";
		wait for Clk_period;
		Addr <=  "00101101111100";
		Trees_din <= x"ffda2ead";
		wait for Clk_period;
		Addr <=  "00101101111101";
		Trees_din <= x"1b004304";
		wait for Clk_period;
		Addr <=  "00101101111110";
		Trees_din <= x"ff952ead";
		wait for Clk_period;
		Addr <=  "00101101111111";
		Trees_din <= x"00242ead";
		wait for Clk_period;
		Addr <=  "00101110000000";
		Trees_din <= x"02ffbf2c";
		wait for Clk_period;
		Addr <=  "00101110000001";
		Trees_din <= x"06f68b10";
		wait for Clk_period;
		Addr <=  "00101110000010";
		Trees_din <= x"1c002704";
		wait for Clk_period;
		Addr <=  "00101110000011";
		Trees_din <= x"ffe22ead";
		wait for Clk_period;
		Addr <=  "00101110000100";
		Trees_din <= x"010fd308";
		wait for Clk_period;
		Addr <=  "00101110000101";
		Trees_din <= x"18004e04";
		wait for Clk_period;
		Addr <=  "00101110000110";
		Trees_din <= x"00852ead";
		wait for Clk_period;
		Addr <=  "00101110000111";
		Trees_din <= x"00052ead";
		wait for Clk_period;
		Addr <=  "00101110001000";
		Trees_din <= x"fffa2ead";
		wait for Clk_period;
		Addr <=  "00101110001001";
		Trees_din <= x"0f02af10";
		wait for Clk_period;
		Addr <=  "00101110001010";
		Trees_din <= x"12033908";
		wait for Clk_period;
		Addr <=  "00101110001011";
		Trees_din <= x"14014304";
		wait for Clk_period;
		Addr <=  "00101110001100";
		Trees_din <= x"00042ead";
		wait for Clk_period;
		Addr <=  "00101110001101";
		Trees_din <= x"00712ead";
		wait for Clk_period;
		Addr <=  "00101110001110";
		Trees_din <= x"09005204";
		wait for Clk_period;
		Addr <=  "00101110001111";
		Trees_din <= x"001b2ead";
		wait for Clk_period;
		Addr <=  "00101110010000";
		Trees_din <= x"ff9c2ead";
		wait for Clk_period;
		Addr <=  "00101110010001";
		Trees_din <= x"11028608";
		wait for Clk_period;
		Addr <=  "00101110010010";
		Trees_din <= x"17000104";
		wait for Clk_period;
		Addr <=  "00101110010011";
		Trees_din <= x"ffe72ead";
		wait for Clk_period;
		Addr <=  "00101110010100";
		Trees_din <= x"ff552ead";
		wait for Clk_period;
		Addr <=  "00101110010101";
		Trees_din <= x"00382ead";
		wait for Clk_period;
		Addr <=  "00101110010110";
		Trees_din <= x"13f83c0c";
		wait for Clk_period;
		Addr <=  "00101110010111";
		Trees_din <= x"19009b08";
		wait for Clk_period;
		Addr <=  "00101110011000";
		Trees_din <= x"0c004604";
		wait for Clk_period;
		Addr <=  "00101110011001";
		Trees_din <= x"fffc2ead";
		wait for Clk_period;
		Addr <=  "00101110011010";
		Trees_din <= x"ff6d2ead";
		wait for Clk_period;
		Addr <=  "00101110011011";
		Trees_din <= x"00432ead";
		wait for Clk_period;
		Addr <=  "00101110011100";
		Trees_din <= x"13f8f710";
		wait for Clk_period;
		Addr <=  "00101110011101";
		Trees_din <= x"06f67408";
		wait for Clk_period;
		Addr <=  "00101110011110";
		Trees_din <= x"05fbe004";
		wait for Clk_period;
		Addr <=  "00101110011111";
		Trees_din <= x"00822ead";
		wait for Clk_period;
		Addr <=  "00101110100000";
		Trees_din <= x"fff62ead";
		wait for Clk_period;
		Addr <=  "00101110100001";
		Trees_din <= x"0109bf04";
		wait for Clk_period;
		Addr <=  "00101110100010";
		Trees_din <= x"00312ead";
		wait for Clk_period;
		Addr <=  "00101110100011";
		Trees_din <= x"ffab2ead";
		wait for Clk_period;
		Addr <=  "00101110100100";
		Trees_din <= x"13019608";
		wait for Clk_period;
		Addr <=  "00101110100101";
		Trees_din <= x"06fb4b04";
		wait for Clk_period;
		Addr <=  "00101110100110";
		Trees_din <= x"fff52ead";
		wait for Clk_period;
		Addr <=  "00101110100111";
		Trees_din <= x"00332ead";
		wait for Clk_period;
		Addr <=  "00101110101000";
		Trees_din <= x"17011904";
		wait for Clk_period;
		Addr <=  "00101110101001";
		Trees_din <= x"00032ead";
		wait for Clk_period;
		Addr <=  "00101110101010";
		Trees_din <= x"006f2ead";
		wait for Clk_period;
		Addr <=  "00101110101011";
		Trees_din <= x"000fd344";
		wait for Clk_period;
		Addr <=  "00101110101100";
		Trees_din <= x"09005d38";
		wait for Clk_period;
		Addr <=  "00101110101101";
		Trees_din <= x"020c6020";
		wait for Clk_period;
		Addr <=  "00101110101110";
		Trees_din <= x"06f73010";
		wait for Clk_period;
		Addr <=  "00101110101111";
		Trees_din <= x"13f88908";
		wait for Clk_period;
		Addr <=  "00101110110000";
		Trees_din <= x"0a026704";
		wait for Clk_period;
		Addr <=  "00101110110001";
		Trees_din <= x"000d2fe1";
		wait for Clk_period;
		Addr <=  "00101110110010";
		Trees_din <= x"ff7a2fe1";
		wait for Clk_period;
		Addr <=  "00101110110011";
		Trees_din <= x"13f8b404";
		wait for Clk_period;
		Addr <=  "00101110110100";
		Trees_din <= x"006d2fe1";
		wait for Clk_period;
		Addr <=  "00101110110101";
		Trees_din <= x"00062fe1";
		wait for Clk_period;
		Addr <=  "00101110110110";
		Trees_din <= x"08019908";
		wait for Clk_period;
		Addr <=  "00101110110111";
		Trees_din <= x"15009a04";
		wait for Clk_period;
		Addr <=  "00101110111000";
		Trees_din <= x"fff02fe1";
		wait for Clk_period;
		Addr <=  "00101110111001";
		Trees_din <= x"ff9b2fe1";
		wait for Clk_period;
		Addr <=  "00101110111010";
		Trees_din <= x"0a02b204";
		wait for Clk_period;
		Addr <=  "00101110111011";
		Trees_din <= x"00312fe1";
		wait for Clk_period;
		Addr <=  "00101110111100";
		Trees_din <= x"ffa92fe1";
		wait for Clk_period;
		Addr <=  "00101110111101";
		Trees_din <= x"06f5b40c";
		wait for Clk_period;
		Addr <=  "00101110111110";
		Trees_din <= x"000e9004";
		wait for Clk_period;
		Addr <=  "00101110111111";
		Trees_din <= x"ff742fe1";
		wait for Clk_period;
		Addr <=  "00101111000000";
		Trees_din <= x"06f46e04";
		wait for Clk_period;
		Addr <=  "00101111000001";
		Trees_din <= x"004a2fe1";
		wait for Clk_period;
		Addr <=  "00101111000010";
		Trees_din <= x"ffa52fe1";
		wait for Clk_period;
		Addr <=  "00101111000011";
		Trees_din <= x"18004308";
		wait for Clk_period;
		Addr <=  "00101111000100";
		Trees_din <= x"1c003204";
		wait for Clk_period;
		Addr <=  "00101111000101";
		Trees_din <= x"fff52fe1";
		wait for Clk_period;
		Addr <=  "00101111000110";
		Trees_din <= x"00882fe1";
		wait for Clk_period;
		Addr <=  "00101111000111";
		Trees_din <= x"ffa42fe1";
		wait for Clk_period;
		Addr <=  "00101111001000";
		Trees_din <= x"04ffda08";
		wait for Clk_period;
		Addr <=  "00101111001001";
		Trees_din <= x"12010b04";
		wait for Clk_period;
		Addr <=  "00101111001010";
		Trees_din <= x"000f2fe1";
		wait for Clk_period;
		Addr <=  "00101111001011";
		Trees_din <= x"007f2fe1";
		wait for Clk_period;
		Addr <=  "00101111001100";
		Trees_din <= x"ffe22fe1";
		wait for Clk_period;
		Addr <=  "00101111001101";
		Trees_din <= x"0afb1130";
		wait for Clk_period;
		Addr <=  "00101111001110";
		Trees_din <= x"1a00c518";
		wait for Clk_period;
		Addr <=  "00101111001111";
		Trees_din <= x"0011920c";
		wait for Clk_period;
		Addr <=  "00101111010000";
		Trees_din <= x"05fb5608";
		wait for Clk_period;
		Addr <=  "00101111010001";
		Trees_din <= x"04fa6f04";
		wait for Clk_period;
		Addr <=  "00101111010010";
		Trees_din <= x"ff682fe1";
		wait for Clk_period;
		Addr <=  "00101111010011";
		Trees_din <= x"fffd2fe1";
		wait for Clk_period;
		Addr <=  "00101111010100";
		Trees_din <= x"00542fe1";
		wait for Clk_period;
		Addr <=  "00101111010101";
		Trees_din <= x"02039104";
		wait for Clk_period;
		Addr <=  "00101111010110";
		Trees_din <= x"007a2fe1";
		wait for Clk_period;
		Addr <=  "00101111010111";
		Trees_din <= x"0f014a04";
		wait for Clk_period;
		Addr <=  "00101111011000";
		Trees_din <= x"00452fe1";
		wait for Clk_period;
		Addr <=  "00101111011001";
		Trees_din <= x"ffc72fe1";
		wait for Clk_period;
		Addr <=  "00101111011010";
		Trees_din <= x"18003b08";
		wait for Clk_period;
		Addr <=  "00101111011011";
		Trees_din <= x"0d010904";
		wait for Clk_period;
		Addr <=  "00101111011100";
		Trees_din <= x"ffd42fe1";
		wait for Clk_period;
		Addr <=  "00101111011101";
		Trees_din <= x"007a2fe1";
		wait for Clk_period;
		Addr <=  "00101111011110";
		Trees_din <= x"11011308";
		wait for Clk_period;
		Addr <=  "00101111011111";
		Trees_din <= x"10042304";
		wait for Clk_period;
		Addr <=  "00101111100000";
		Trees_din <= x"ffe72fe1";
		wait for Clk_period;
		Addr <=  "00101111100001";
		Trees_din <= x"00562fe1";
		wait for Clk_period;
		Addr <=  "00101111100010";
		Trees_din <= x"15009704";
		wait for Clk_period;
		Addr <=  "00101111100011";
		Trees_din <= x"ffed2fe1";
		wait for Clk_period;
		Addr <=  "00101111100100";
		Trees_din <= x"ff632fe1";
		wait for Clk_period;
		Addr <=  "00101111100101";
		Trees_din <= x"0afb2608";
		wait for Clk_period;
		Addr <=  "00101111100110";
		Trees_din <= x"08009604";
		wait for Clk_period;
		Addr <=  "00101111100111";
		Trees_din <= x"002c2fe1";
		wait for Clk_period;
		Addr <=  "00101111101000";
		Trees_din <= x"00982fe1";
		wait for Clk_period;
		Addr <=  "00101111101001";
		Trees_din <= x"010b3210";
		wait for Clk_period;
		Addr <=  "00101111101010";
		Trees_din <= x"08015708";
		wait for Clk_period;
		Addr <=  "00101111101011";
		Trees_din <= x"0e043204";
		wait for Clk_period;
		Addr <=  "00101111101100";
		Trees_din <= x"006e2fe1";
		wait for Clk_period;
		Addr <=  "00101111101101";
		Trees_din <= x"ffe32fe1";
		wait for Clk_period;
		Addr <=  "00101111101110";
		Trees_din <= x"1900a504";
		wait for Clk_period;
		Addr <=  "00101111101111";
		Trees_din <= x"ffeb2fe1";
		wait for Clk_period;
		Addr <=  "00101111110000";
		Trees_din <= x"00692fe1";
		wait for Clk_period;
		Addr <=  "00101111110001";
		Trees_din <= x"05f9fc08";
		wait for Clk_period;
		Addr <=  "00101111110010";
		Trees_din <= x"0c024504";
		wait for Clk_period;
		Addr <=  "00101111110011";
		Trees_din <= x"00492fe1";
		wait for Clk_period;
		Addr <=  "00101111110100";
		Trees_din <= x"ffe02fe1";
		wait for Clk_period;
		Addr <=  "00101111110101";
		Trees_din <= x"15008504";
		wait for Clk_period;
		Addr <=  "00101111110110";
		Trees_din <= x"006b2fe1";
		wait for Clk_period;
		Addr <=  "00101111110111";
		Trees_din <= x"ffc62fe1";
		wait for Clk_period;
		Addr <=  "00101111111000";
		Trees_din <= x"000b1e4c";
		wait for Clk_period;
		Addr <=  "00101111111001";
		Trees_din <= x"18003d24";
		wait for Clk_period;
		Addr <=  "00101111111010";
		Trees_din <= x"1c002f18";
		wait for Clk_period;
		Addr <=  "00101111111011";
		Trees_din <= x"1103d610";
		wait for Clk_period;
		Addr <=  "00101111111100";
		Trees_din <= x"0e00ea08";
		wait for Clk_period;
		Addr <=  "00101111111101";
		Trees_din <= x"04fbe704";
		wait for Clk_period;
		Addr <=  "00101111111110";
		Trees_din <= x"005d312d";
		wait for Clk_period;
		Addr <=  "00101111111111";
		Trees_din <= x"ff94312d";
		wait for Clk_period;
		Addr <=  "00110000000000";
		Trees_din <= x"0bf95304";
		wait for Clk_period;
		Addr <=  "00110000000001";
		Trees_din <= x"ffcc312d";
		wait for Clk_period;
		Addr <=  "00110000000010";
		Trees_din <= x"0045312d";
		wait for Clk_period;
		Addr <=  "00110000000011";
		Trees_din <= x"00050804";
		wait for Clk_period;
		Addr <=  "00110000000100";
		Trees_din <= x"fffa312d";
		wait for Clk_period;
		Addr <=  "00110000000101";
		Trees_din <= x"ff73312d";
		wait for Clk_period;
		Addr <=  "00110000000110";
		Trees_din <= x"1a00d508";
		wait for Clk_period;
		Addr <=  "00110000000111";
		Trees_din <= x"14034004";
		wait for Clk_period;
		Addr <=  "00110000001000";
		Trees_din <= x"ffbe312d";
		wait for Clk_period;
		Addr <=  "00110000001001";
		Trees_din <= x"002b312d";
		wait for Clk_period;
		Addr <=  "00110000001010";
		Trees_din <= x"ff71312d";
		wait for Clk_period;
		Addr <=  "00110000001011";
		Trees_din <= x"1b003308";
		wait for Clk_period;
		Addr <=  "00110000001100";
		Trees_din <= x"14026e04";
		wait for Clk_period;
		Addr <=  "00110000001101";
		Trees_din <= x"008b312d";
		wait for Clk_period;
		Addr <=  "00110000001110";
		Trees_din <= x"ffef312d";
		wait for Clk_period;
		Addr <=  "00110000001111";
		Trees_din <= x"17018e10";
		wait for Clk_period;
		Addr <=  "00110000010000";
		Trees_din <= x"0b056f08";
		wait for Clk_period;
		Addr <=  "00110000010001";
		Trees_din <= x"12028704";
		wait for Clk_period;
		Addr <=  "00110000010010";
		Trees_din <= x"ffc4312d";
		wait for Clk_period;
		Addr <=  "00110000010011";
		Trees_din <= x"000b312d";
		wait for Clk_period;
		Addr <=  "00110000010100";
		Trees_din <= x"07005804";
		wait for Clk_period;
		Addr <=  "00110000010101";
		Trees_din <= x"0083312d";
		wait for Clk_period;
		Addr <=  "00110000010110";
		Trees_din <= x"ffa2312d";
		wait for Clk_period;
		Addr <=  "00110000010111";
		Trees_din <= x"0d01e508";
		wait for Clk_period;
		Addr <=  "00110000011000";
		Trees_din <= x"07005604";
		wait for Clk_period;
		Addr <=  "00110000011001";
		Trees_din <= x"004c312d";
		wait for Clk_period;
		Addr <=  "00110000011010";
		Trees_din <= x"ffdf312d";
		wait for Clk_period;
		Addr <=  "00110000011011";
		Trees_din <= x"1603f704";
		wait for Clk_period;
		Addr <=  "00110000011100";
		Trees_din <= x"0069312d";
		wait for Clk_period;
		Addr <=  "00110000011101";
		Trees_din <= x"ffc4312d";
		wait for Clk_period;
		Addr <=  "00110000011110";
		Trees_din <= x"0105aa24";
		wait for Clk_period;
		Addr <=  "00110000011111";
		Trees_din <= x"1b002f04";
		wait for Clk_period;
		Addr <=  "00110000100000";
		Trees_din <= x"0080312d";
		wait for Clk_period;
		Addr <=  "00110000100001";
		Trees_din <= x"1e006110";
		wait for Clk_period;
		Addr <=  "00110000100010";
		Trees_din <= x"05fcab08";
		wait for Clk_period;
		Addr <=  "00110000100011";
		Trees_din <= x"1400fd04";
		wait for Clk_period;
		Addr <=  "00110000100100";
		Trees_din <= x"fffa312d";
		wait for Clk_period;
		Addr <=  "00110000100101";
		Trees_din <= x"0069312d";
		wait for Clk_period;
		Addr <=  "00110000100110";
		Trees_din <= x"16037804";
		wait for Clk_period;
		Addr <=  "00110000100111";
		Trees_din <= x"ff9d312d";
		wait for Clk_period;
		Addr <=  "00110000101000";
		Trees_din <= x"0042312d";
		wait for Clk_period;
		Addr <=  "00110000101001";
		Trees_din <= x"08003408";
		wait for Clk_period;
		Addr <=  "00110000101010";
		Trees_din <= x"0d01d504";
		wait for Clk_period;
		Addr <=  "00110000101011";
		Trees_din <= x"0050312d";
		wait for Clk_period;
		Addr <=  "00110000101100";
		Trees_din <= x"ffc2312d";
		wait for Clk_period;
		Addr <=  "00110000101101";
		Trees_din <= x"07005804";
		wait for Clk_period;
		Addr <=  "00110000101110";
		Trees_din <= x"001a312d";
		wait for Clk_period;
		Addr <=  "00110000101111";
		Trees_din <= x"0074312d";
		wait for Clk_period;
		Addr <=  "00110000110000";
		Trees_din <= x"02ffe318";
		wait for Clk_period;
		Addr <=  "00110000110001";
		Trees_din <= x"13ffb70c";
		wait for Clk_period;
		Addr <=  "00110000110010";
		Trees_din <= x"000f3608";
		wait for Clk_period;
		Addr <=  "00110000110011";
		Trees_din <= x"03fa9f04";
		wait for Clk_period;
		Addr <=  "00110000110100";
		Trees_din <= x"ffb4312d";
		wait for Clk_period;
		Addr <=  "00110000110101";
		Trees_din <= x"0064312d";
		wait for Clk_period;
		Addr <=  "00110000110110";
		Trees_din <= x"0083312d";
		wait for Clk_period;
		Addr <=  "00110000110111";
		Trees_din <= x"09005404";
		wait for Clk_period;
		Addr <=  "00110000111000";
		Trees_din <= x"0056312d";
		wait for Clk_period;
		Addr <=  "00110000111001";
		Trees_din <= x"15009904";
		wait for Clk_period;
		Addr <=  "00110000111010";
		Trees_din <= x"ff7a312d";
		wait for Clk_period;
		Addr <=  "00110000111011";
		Trees_din <= x"0008312d";
		wait for Clk_period;
		Addr <=  "00110000111100";
		Trees_din <= x"05f7e710";
		wait for Clk_period;
		Addr <=  "00110000111101";
		Trees_din <= x"0a031a08";
		wait for Clk_period;
		Addr <=  "00110000111110";
		Trees_din <= x"1500a404";
		wait for Clk_period;
		Addr <=  "00110000111111";
		Trees_din <= x"0053312d";
		wait for Clk_period;
		Addr <=  "00110001000000";
		Trees_din <= x"ffe4312d";
		wait for Clk_period;
		Addr <=  "00110001000001";
		Trees_din <= x"0205a104";
		wait for Clk_period;
		Addr <=  "00110001000010";
		Trees_din <= x"fff1312d";
		wait for Clk_period;
		Addr <=  "00110001000011";
		Trees_din <= x"ff98312d";
		wait for Clk_period;
		Addr <=  "00110001000100";
		Trees_din <= x"07005b08";
		wait for Clk_period;
		Addr <=  "00110001000101";
		Trees_din <= x"07005a04";
		wait for Clk_period;
		Addr <=  "00110001000110";
		Trees_din <= x"fff6312d";
		wait for Clk_period;
		Addr <=  "00110001000111";
		Trees_din <= x"0067312d";
		wait for Clk_period;
		Addr <=  "00110001001000";
		Trees_din <= x"10fa4504";
		wait for Clk_period;
		Addr <=  "00110001001001";
		Trees_din <= x"0062312d";
		wait for Clk_period;
		Addr <=  "00110001001010";
		Trees_din <= x"ffa3312d";
		wait for Clk_period;
		Addr <=  "00110001001011";
		Trees_din <= x"000fd350";
		wait for Clk_period;
		Addr <=  "00110001001100";
		Trees_din <= x"11fe7224";
		wait for Clk_period;
		Addr <=  "00110001001101";
		Trees_din <= x"1c003510";
		wait for Clk_period;
		Addr <=  "00110001001110";
		Trees_din <= x"1603d10c";
		wait for Clk_period;
		Addr <=  "00110001001111";
		Trees_din <= x"0f000f04";
		wait for Clk_period;
		Addr <=  "00110001010000";
		Trees_din <= x"000c3259";
		wait for Clk_period;
		Addr <=  "00110001010001";
		Trees_din <= x"0101d104";
		wait for Clk_period;
		Addr <=  "00110001010010";
		Trees_din <= x"ffd23259";
		wait for Clk_period;
		Addr <=  "00110001010011";
		Trees_din <= x"ff623259";
		wait for Clk_period;
		Addr <=  "00110001010100";
		Trees_din <= x"00363259";
		wait for Clk_period;
		Addr <=  "00110001010101";
		Trees_din <= x"1b003504";
		wait for Clk_period;
		Addr <=  "00110001010110";
		Trees_din <= x"00773259";
		wait for Clk_period;
		Addr <=  "00110001010111";
		Trees_din <= x"13ffd008";
		wait for Clk_period;
		Addr <=  "00110001011000";
		Trees_din <= x"14016004";
		wait for Clk_period;
		Addr <=  "00110001011001";
		Trees_din <= x"00103259";
		wait for Clk_period;
		Addr <=  "00110001011010";
		Trees_din <= x"ff823259";
		wait for Clk_period;
		Addr <=  "00110001011011";
		Trees_din <= x"1b003e04";
		wait for Clk_period;
		Addr <=  "00110001011100";
		Trees_din <= x"ffda3259";
		wait for Clk_period;
		Addr <=  "00110001011101";
		Trees_din <= x"00653259";
		wait for Clk_period;
		Addr <=  "00110001011110";
		Trees_din <= x"0a044c20";
		wait for Clk_period;
		Addr <=  "00110001011111";
		Trees_din <= x"19008710";
		wait for Clk_period;
		Addr <=  "00110001100000";
		Trees_din <= x"05fb8408";
		wait for Clk_period;
		Addr <=  "00110001100001";
		Trees_din <= x"11ff2e04";
		wait for Clk_period;
		Addr <=  "00110001100010";
		Trees_din <= x"00353259";
		wait for Clk_period;
		Addr <=  "00110001100011";
		Trees_din <= x"ff923259";
		wait for Clk_period;
		Addr <=  "00110001100100";
		Trees_din <= x"08002604";
		wait for Clk_period;
		Addr <=  "00110001100101";
		Trees_din <= x"ffbd3259";
		wait for Clk_period;
		Addr <=  "00110001100110";
		Trees_din <= x"002a3259";
		wait for Clk_period;
		Addr <=  "00110001100111";
		Trees_din <= x"0bfa4108";
		wait for Clk_period;
		Addr <=  "00110001101000";
		Trees_din <= x"08001504";
		wait for Clk_period;
		Addr <=  "00110001101001";
		Trees_din <= x"00503259";
		wait for Clk_period;
		Addr <=  "00110001101010";
		Trees_din <= x"ffce3259";
		wait for Clk_period;
		Addr <=  "00110001101011";
		Trees_din <= x"1e005a04";
		wait for Clk_period;
		Addr <=  "00110001101100";
		Trees_din <= x"ffd83259";
		wait for Clk_period;
		Addr <=  "00110001101101";
		Trees_din <= x"001b3259";
		wait for Clk_period;
		Addr <=  "00110001101110";
		Trees_din <= x"11ff0608";
		wait for Clk_period;
		Addr <=  "00110001101111";
		Trees_din <= x"04faa904";
		wait for Clk_period;
		Addr <=  "00110001110000";
		Trees_din <= x"005a3259";
		wait for Clk_period;
		Addr <=  "00110001110001";
		Trees_din <= x"ffc43259";
		wait for Clk_period;
		Addr <=  "00110001110010";
		Trees_din <= x"008b3259";
		wait for Clk_period;
		Addr <=  "00110001110011";
		Trees_din <= x"0afb1124";
		wait for Clk_period;
		Addr <=  "00110001110100";
		Trees_din <= x"00119210";
		wait for Clk_period;
		Addr <=  "00110001110101";
		Trees_din <= x"0e007004";
		wait for Clk_period;
		Addr <=  "00110001110110";
		Trees_din <= x"00323259";
		wait for Clk_period;
		Addr <=  "00110001110111";
		Trees_din <= x"1500a408";
		wait for Clk_period;
		Addr <=  "00110001111000";
		Trees_din <= x"02079804";
		wait for Clk_period;
		Addr <=  "00110001111001";
		Trees_din <= x"ff703259";
		wait for Clk_period;
		Addr <=  "00110001111010";
		Trees_din <= x"fff03259";
		wait for Clk_period;
		Addr <=  "00110001111011";
		Trees_din <= x"00133259";
		wait for Clk_period;
		Addr <=  "00110001111100";
		Trees_din <= x"09005004";
		wait for Clk_period;
		Addr <=  "00110001111101";
		Trees_din <= x"006f3259";
		wait for Clk_period;
		Addr <=  "00110001111110";
		Trees_din <= x"1a00c708";
		wait for Clk_period;
		Addr <=  "00110001111111";
		Trees_din <= x"02039104";
		wait for Clk_period;
		Addr <=  "00110010000000";
		Trees_din <= x"00753259";
		wait for Clk_period;
		Addr <=  "00110010000001";
		Trees_din <= x"00033259";
		wait for Clk_period;
		Addr <=  "00110010000010";
		Trees_din <= x"1c003104";
		wait for Clk_period;
		Addr <=  "00110010000011";
		Trees_din <= x"00193259";
		wait for Clk_period;
		Addr <=  "00110010000100";
		Trees_din <= x"ff893259";
		wait for Clk_period;
		Addr <=  "00110010000101";
		Trees_din <= x"0afb2604";
		wait for Clk_period;
		Addr <=  "00110010000110";
		Trees_din <= x"00843259";
		wait for Clk_period;
		Addr <=  "00110010000111";
		Trees_din <= x"06f71110";
		wait for Clk_period;
		Addr <=  "00110010001000";
		Trees_din <= x"0afccc08";
		wait for Clk_period;
		Addr <=  "00110010001001";
		Trees_din <= x"05f9ce04";
		wait for Clk_period;
		Addr <=  "00110010001010";
		Trees_din <= x"001f3259";
		wait for Clk_period;
		Addr <=  "00110010001011";
		Trees_din <= x"ffaa3259";
		wait for Clk_period;
		Addr <=  "00110010001100";
		Trees_din <= x"1c002d04";
		wait for Clk_period;
		Addr <=  "00110010001101";
		Trees_din <= x"00603259";
		wait for Clk_period;
		Addr <=  "00110010001110";
		Trees_din <= x"fffe3259";
		wait for Clk_period;
		Addr <=  "00110010001111";
		Trees_din <= x"0eff2d08";
		wait for Clk_period;
		Addr <=  "00110010010000";
		Trees_din <= x"0d030d04";
		wait for Clk_period;
		Addr <=  "00110010010001";
		Trees_din <= x"002d3259";
		wait for Clk_period;
		Addr <=  "00110010010010";
		Trees_din <= x"ffa13259";
		wait for Clk_period;
		Addr <=  "00110010010011";
		Trees_din <= x"02075104";
		wait for Clk_period;
		Addr <=  "00110010010100";
		Trees_din <= x"006e3259";
		wait for Clk_period;
		Addr <=  "00110010010101";
		Trees_din <= x"ffe73259";
		wait for Clk_period;
		Addr <=  "00110010010110";
		Trees_din <= x"0111ec74";
		wait for Clk_period;
		Addr <=  "00110010010111";
		Trees_din <= x"03f78338";
		wait for Clk_period;
		Addr <=  "00110010011000";
		Trees_din <= x"0c00b718";
		wait for Clk_period;
		Addr <=  "00110010011001";
		Trees_din <= x"1201d60c";
		wait for Clk_period;
		Addr <=  "00110010011010";
		Trees_din <= x"13ffc508";
		wait for Clk_period;
		Addr <=  "00110010011011";
		Trees_din <= x"07005b04";
		wait for Clk_period;
		Addr <=  "00110010011100";
		Trees_din <= x"006633a5";
		wait for Clk_period;
		Addr <=  "00110010011101";
		Trees_din <= x"fff333a5";
		wait for Clk_period;
		Addr <=  "00110010011110";
		Trees_din <= x"ffbe33a5";
		wait for Clk_period;
		Addr <=  "00110010011111";
		Trees_din <= x"04f90008";
		wait for Clk_period;
		Addr <=  "00110010100000";
		Trees_din <= x"1a00cc04";
		wait for Clk_period;
		Addr <=  "00110010100001";
		Trees_din <= x"ffc533a5";
		wait for Clk_period;
		Addr <=  "00110010100010";
		Trees_din <= x"004a33a5";
		wait for Clk_period;
		Addr <=  "00110010100011";
		Trees_din <= x"ff6133a5";
		wait for Clk_period;
		Addr <=  "00110010100100";
		Trees_din <= x"02094410";
		wait for Clk_period;
		Addr <=  "00110010100101";
		Trees_din <= x"07005808";
		wait for Clk_period;
		Addr <=  "00110010100110";
		Trees_din <= x"0800af04";
		wait for Clk_period;
		Addr <=  "00110010100111";
		Trees_din <= x"000933a5";
		wait for Clk_period;
		Addr <=  "00110010101000";
		Trees_din <= x"007e33a5";
		wait for Clk_period;
		Addr <=  "00110010101001";
		Trees_din <= x"17000204";
		wait for Clk_period;
		Addr <=  "00110010101010";
		Trees_din <= x"006033a5";
		wait for Clk_period;
		Addr <=  "00110010101011";
		Trees_din <= x"ffde33a5";
		wait for Clk_period;
		Addr <=  "00110010101100";
		Trees_din <= x"010e3108";
		wait for Clk_period;
		Addr <=  "00110010101101";
		Trees_din <= x"000f0704";
		wait for Clk_period;
		Addr <=  "00110010101110";
		Trees_din <= x"ffaf33a5";
		wait for Clk_period;
		Addr <=  "00110010101111";
		Trees_din <= x"002533a5";
		wait for Clk_period;
		Addr <=  "00110010110000";
		Trees_din <= x"0afb6204";
		wait for Clk_period;
		Addr <=  "00110010110001";
		Trees_din <= x"fff633a5";
		wait for Clk_period;
		Addr <=  "00110010110010";
		Trees_din <= x"ff8733a5";
		wait for Clk_period;
		Addr <=  "00110010110011";
		Trees_din <= x"0c038320";
		wait for Clk_period;
		Addr <=  "00110010110100";
		Trees_din <= x"0af7cc10";
		wait for Clk_period;
		Addr <=  "00110010110101";
		Trees_din <= x"0102a908";
		wait for Clk_period;
		Addr <=  "00110010110110";
		Trees_din <= x"01009804";
		wait for Clk_period;
		Addr <=  "00110010110111";
		Trees_din <= x"fffe33a5";
		wait for Clk_period;
		Addr <=  "00110010111000";
		Trees_din <= x"007133a5";
		wait for Clk_period;
		Addr <=  "00110010111001";
		Trees_din <= x"08003004";
		wait for Clk_period;
		Addr <=  "00110010111010";
		Trees_din <= x"fff833a5";
		wait for Clk_period;
		Addr <=  "00110010111011";
		Trees_din <= x"ff7c33a5";
		wait for Clk_period;
		Addr <=  "00110010111100";
		Trees_din <= x"11021b08";
		wait for Clk_period;
		Addr <=  "00110010111101";
		Trees_din <= x"05ffdf04";
		wait for Clk_period;
		Addr <=  "00110010111110";
		Trees_din <= x"002033a5";
		wait for Clk_period;
		Addr <=  "00110010111111";
		Trees_din <= x"ffaa33a5";
		wait for Clk_period;
		Addr <=  "00110011000000";
		Trees_din <= x"07005a04";
		wait for Clk_period;
		Addr <=  "00110011000001";
		Trees_din <= x"ffed33a5";
		wait for Clk_period;
		Addr <=  "00110011000010";
		Trees_din <= x"002233a5";
		wait for Clk_period;
		Addr <=  "00110011000011";
		Trees_din <= x"0108a410";
		wait for Clk_period;
		Addr <=  "00110011000100";
		Trees_din <= x"06f4ea08";
		wait for Clk_period;
		Addr <=  "00110011000101";
		Trees_din <= x"0afaec04";
		wait for Clk_period;
		Addr <=  "00110011000110";
		Trees_din <= x"006b33a5";
		wait for Clk_period;
		Addr <=  "00110011000111";
		Trees_din <= x"000d33a5";
		wait for Clk_period;
		Addr <=  "00110011001000";
		Trees_din <= x"19009f04";
		wait for Clk_period;
		Addr <=  "00110011001001";
		Trees_din <= x"ffbb33a5";
		wait for Clk_period;
		Addr <=  "00110011001010";
		Trees_din <= x"003c33a5";
		wait for Clk_period;
		Addr <=  "00110011001011";
		Trees_din <= x"02ffc504";
		wait for Clk_period;
		Addr <=  "00110011001100";
		Trees_din <= x"002433a5";
		wait for Clk_period;
		Addr <=  "00110011001101";
		Trees_din <= x"1500a004";
		wait for Clk_period;
		Addr <=  "00110011001110";
		Trees_din <= x"ff7533a5";
		wait for Clk_period;
		Addr <=  "00110011001111";
		Trees_din <= x"ffe733a5";
		wait for Clk_period;
		Addr <=  "00110011010000";
		Trees_din <= x"14006604";
		wait for Clk_period;
		Addr <=  "00110011010001";
		Trees_din <= x"ff8b33a5";
		wait for Clk_period;
		Addr <=  "00110011010010";
		Trees_din <= x"06f4f214";
		wait for Clk_period;
		Addr <=  "00110011010011";
		Trees_din <= x"1d004e0c";
		wait for Clk_period;
		Addr <=  "00110011010100";
		Trees_din <= x"0c00d704";
		wait for Clk_period;
		Addr <=  "00110011010101";
		Trees_din <= x"000133a5";
		wait for Clk_period;
		Addr <=  "00110011010110";
		Trees_din <= x"11012204";
		wait for Clk_period;
		Addr <=  "00110011010111";
		Trees_din <= x"ffe133a5";
		wait for Clk_period;
		Addr <=  "00110011011000";
		Trees_din <= x"ff8133a5";
		wait for Clk_period;
		Addr <=  "00110011011001";
		Trees_din <= x"11027c04";
		wait for Clk_period;
		Addr <=  "00110011011010";
		Trees_din <= x"ffe933a5";
		wait for Clk_period;
		Addr <=  "00110011011011";
		Trees_din <= x"005f33a5";
		wait for Clk_period;
		Addr <=  "00110011011100";
		Trees_din <= x"06f57f0c";
		wait for Clk_period;
		Addr <=  "00110011011101";
		Trees_din <= x"1d004004";
		wait for Clk_period;
		Addr <=  "00110011011110";
		Trees_din <= x"fff033a5";
		wait for Clk_period;
		Addr <=  "00110011011111";
		Trees_din <= x"1c003704";
		wait for Clk_period;
		Addr <=  "00110011100000";
		Trees_din <= x"00af33a5";
		wait for Clk_period;
		Addr <=  "00110011100001";
		Trees_din <= x"002933a5";
		wait for Clk_period;
		Addr <=  "00110011100010";
		Trees_din <= x"1401ad08";
		wait for Clk_period;
		Addr <=  "00110011100011";
		Trees_din <= x"0011ff04";
		wait for Clk_period;
		Addr <=  "00110011100100";
		Trees_din <= x"fff433a5";
		wait for Clk_period;
		Addr <=  "00110011100101";
		Trees_din <= x"005b33a5";
		wait for Clk_period;
		Addr <=  "00110011100110";
		Trees_din <= x"0f02dd04";
		wait for Clk_period;
		Addr <=  "00110011100111";
		Trees_din <= x"ff8933a5";
		wait for Clk_period;
		Addr <=  "00110011101000";
		Trees_din <= x"000c33a5";
		wait for Clk_period;
		Addr <=  "00110011101001";
		Trees_din <= x"0003aa24";
		wait for Clk_period;
		Addr <=  "00110011101010";
		Trees_din <= x"0bf94004";
		wait for Clk_period;
		Addr <=  "00110011101011";
		Trees_din <= x"00343491";
		wait for Clk_period;
		Addr <=  "00110011101100";
		Trees_din <= x"09005414";
		wait for Clk_period;
		Addr <=  "00110011101101";
		Trees_din <= x"1e006108";
		wait for Clk_period;
		Addr <=  "00110011101110";
		Trees_din <= x"1f000004";
		wait for Clk_period;
		Addr <=  "00110011101111";
		Trees_din <= x"ff9c3491";
		wait for Clk_period;
		Addr <=  "00110011110000";
		Trees_din <= x"000a3491";
		wait for Clk_period;
		Addr <=  "00110011110001";
		Trees_din <= x"19008604";
		wait for Clk_period;
		Addr <=  "00110011110010";
		Trees_din <= x"ffc43491";
		wait for Clk_period;
		Addr <=  "00110011110011";
		Trees_din <= x"10faaa04";
		wait for Clk_period;
		Addr <=  "00110011110100";
		Trees_din <= x"00643491";
		wait for Clk_period;
		Addr <=  "00110011110101";
		Trees_din <= x"000b3491";
		wait for Clk_period;
		Addr <=  "00110011110110";
		Trees_din <= x"01fd7808";
		wait for Clk_period;
		Addr <=  "00110011110111";
		Trees_din <= x"0f037e04";
		wait for Clk_period;
		Addr <=  "00110011111000";
		Trees_din <= x"ffbc3491";
		wait for Clk_period;
		Addr <=  "00110011111001";
		Trees_din <= x"00323491";
		wait for Clk_period;
		Addr <=  "00110011111010";
		Trees_din <= x"ff803491";
		wait for Clk_period;
		Addr <=  "00110011111011";
		Trees_din <= x"02ffbf2c";
		wait for Clk_period;
		Addr <=  "00110011111100";
		Trees_din <= x"06f68b14";
		wait for Clk_period;
		Addr <=  "00110011111101";
		Trees_din <= x"0d039310";
		wait for Clk_period;
		Addr <=  "00110011111110";
		Trees_din <= x"1e007608";
		wait for Clk_period;
		Addr <=  "00110011111111";
		Trees_din <= x"1c002604";
		wait for Clk_period;
		Addr <=  "00110100000000";
		Trees_din <= x"00093491";
		wait for Clk_period;
		Addr <=  "00110100000001";
		Trees_din <= x"007b3491";
		wait for Clk_period;
		Addr <=  "00110100000010";
		Trees_din <= x"13ff9d04";
		wait for Clk_period;
		Addr <=  "00110100000011";
		Trees_din <= x"ffc13491";
		wait for Clk_period;
		Addr <=  "00110100000100";
		Trees_din <= x"00393491";
		wait for Clk_period;
		Addr <=  "00110100000101";
		Trees_din <= x"ffd63491";
		wait for Clk_period;
		Addr <=  "00110100000110";
		Trees_din <= x"0f003e08";
		wait for Clk_period;
		Addr <=  "00110100000111";
		Trees_din <= x"0b041504";
		wait for Clk_period;
		Addr <=  "00110100001000";
		Trees_din <= x"00723491";
		wait for Clk_period;
		Addr <=  "00110100001001";
		Trees_din <= x"fffd3491";
		wait for Clk_period;
		Addr <=  "00110100001010";
		Trees_din <= x"04022408";
		wait for Clk_period;
		Addr <=  "00110100001011";
		Trees_din <= x"04fd9804";
		wait for Clk_period;
		Addr <=  "00110100001100";
		Trees_din <= x"00053491";
		wait for Clk_period;
		Addr <=  "00110100001101";
		Trees_din <= x"ffa83491";
		wait for Clk_period;
		Addr <=  "00110100001110";
		Trees_din <= x"18004404";
		wait for Clk_period;
		Addr <=  "00110100001111";
		Trees_din <= x"00563491";
		wait for Clk_period;
		Addr <=  "00110100010000";
		Trees_din <= x"00013491";
		wait for Clk_period;
		Addr <=  "00110100010001";
		Trees_din <= x"1006461c";
		wait for Clk_period;
		Addr <=  "00110100010010";
		Trees_din <= x"13f83c0c";
		wait for Clk_period;
		Addr <=  "00110100010011";
		Trees_din <= x"19009b08";
		wait for Clk_period;
		Addr <=  "00110100010100";
		Trees_din <= x"09005304";
		wait for Clk_period;
		Addr <=  "00110100010101";
		Trees_din <= x"ffef3491";
		wait for Clk_period;
		Addr <=  "00110100010110";
		Trees_din <= x"ff803491";
		wait for Clk_period;
		Addr <=  "00110100010111";
		Trees_din <= x"00373491";
		wait for Clk_period;
		Addr <=  "00110100011000";
		Trees_din <= x"13f8f708";
		wait for Clk_period;
		Addr <=  "00110100011001";
		Trees_din <= x"06f67404";
		wait for Clk_period;
		Addr <=  "00110100011010";
		Trees_din <= x"00493491";
		wait for Clk_period;
		Addr <=  "00110100011011";
		Trees_din <= x"ffed3491";
		wait for Clk_period;
		Addr <=  "00110100011100";
		Trees_din <= x"07005b04";
		wait for Clk_period;
		Addr <=  "00110100011101";
		Trees_din <= x"00043491";
		wait for Clk_period;
		Addr <=  "00110100011110";
		Trees_din <= x"ffde3491";
		wait for Clk_period;
		Addr <=  "00110100011111";
		Trees_din <= x"01063004";
		wait for Clk_period;
		Addr <=  "00110100100000";
		Trees_din <= x"00253491";
		wait for Clk_period;
		Addr <=  "00110100100001";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00110100100010";
		Trees_din <= x"ffeb3491";
		wait for Clk_period;
		Addr <=  "00110100100011";
		Trees_din <= x"ff893491";
		wait for Clk_period;
		Addr <=  "00110100100100";
		Trees_din <= x"000b1e2c";
		wait for Clk_period;
		Addr <=  "00110100100101";
		Trees_din <= x"03f85a08";
		wait for Clk_period;
		Addr <=  "00110100100110";
		Trees_din <= x"01060b04";
		wait for Clk_period;
		Addr <=  "00110100100111";
		Trees_din <= x"fffb358d";
		wait for Clk_period;
		Addr <=  "00110100101000";
		Trees_din <= x"ff94358d";
		wait for Clk_period;
		Addr <=  "00110100101001";
		Trees_din <= x"11fed310";
		wait for Clk_period;
		Addr <=  "00110100101010";
		Trees_din <= x"0e00d70c";
		wait for Clk_period;
		Addr <=  "00110100101011";
		Trees_din <= x"0c035a08";
		wait for Clk_period;
		Addr <=  "00110100101100";
		Trees_din <= x"1f000004";
		wait for Clk_period;
		Addr <=  "00110100101101";
		Trees_din <= x"ff8b358d";
		wait for Clk_period;
		Addr <=  "00110100101110";
		Trees_din <= x"000c358d";
		wait for Clk_period;
		Addr <=  "00110100101111";
		Trees_din <= x"0005358d";
		wait for Clk_period;
		Addr <=  "00110100110000";
		Trees_din <= x"002c358d";
		wait for Clk_period;
		Addr <=  "00110100110001";
		Trees_din <= x"0a046710";
		wait for Clk_period;
		Addr <=  "00110100110010";
		Trees_din <= x"0202b808";
		wait for Clk_period;
		Addr <=  "00110100110011";
		Trees_din <= x"09005304";
		wait for Clk_period;
		Addr <=  "00110100110100";
		Trees_din <= x"ffc7358d";
		wait for Clk_period;
		Addr <=  "00110100110101";
		Trees_din <= x"0002358d";
		wait for Clk_period;
		Addr <=  "00110100110110";
		Trees_din <= x"02067004";
		wait for Clk_period;
		Addr <=  "00110100110111";
		Trees_din <= x"0032358d";
		wait for Clk_period;
		Addr <=  "00110100111000";
		Trees_din <= x"ffe7358d";
		wait for Clk_period;
		Addr <=  "00110100111001";
		Trees_din <= x"0066358d";
		wait for Clk_period;
		Addr <=  "00110100111010";
		Trees_din <= x"18003618";
		wait for Clk_period;
		Addr <=  "00110100111011";
		Trees_din <= x"010db60c";
		wait for Clk_period;
		Addr <=  "00110100111100";
		Trees_din <= x"020baf08";
		wait for Clk_period;
		Addr <=  "00110100111101";
		Trees_din <= x"18002e04";
		wait for Clk_period;
		Addr <=  "00110100111110";
		Trees_din <= x"fff8358d";
		wait for Clk_period;
		Addr <=  "00110100111111";
		Trees_din <= x"0094358d";
		wait for Clk_period;
		Addr <=  "00110101000000";
		Trees_din <= x"ffed358d";
		wait for Clk_period;
		Addr <=  "00110101000001";
		Trees_din <= x"00115708";
		wait for Clk_period;
		Addr <=  "00110101000010";
		Trees_din <= x"1c002904";
		wait for Clk_period;
		Addr <=  "00110101000011";
		Trees_din <= x"ff9f358d";
		wait for Clk_period;
		Addr <=  "00110101000100";
		Trees_din <= x"001f358d";
		wait for Clk_period;
		Addr <=  "00110101000101";
		Trees_din <= x"0051358d";
		wait for Clk_period;
		Addr <=  "00110101000110";
		Trees_din <= x"1e005c1c";
		wait for Clk_period;
		Addr <=  "00110101000111";
		Trees_din <= x"0202f30c";
		wait for Clk_period;
		Addr <=  "00110101001000";
		Trees_din <= x"13015208";
		wait for Clk_period;
		Addr <=  "00110101001001";
		Trees_din <= x"1500a104";
		wait for Clk_period;
		Addr <=  "00110101001010";
		Trees_din <= x"0039358d";
		wait for Clk_period;
		Addr <=  "00110101001011";
		Trees_din <= x"ffd1358d";
		wait for Clk_period;
		Addr <=  "00110101001100";
		Trees_din <= x"007f358d";
		wait for Clk_period;
		Addr <=  "00110101001101";
		Trees_din <= x"0f00cf08";
		wait for Clk_period;
		Addr <=  "00110101001110";
		Trees_din <= x"1a00f204";
		wait for Clk_period;
		Addr <=  "00110101001111";
		Trees_din <= x"ff7e358d";
		wait for Clk_period;
		Addr <=  "00110101010000";
		Trees_din <= x"ffe6358d";
		wait for Clk_period;
		Addr <=  "00110101010001";
		Trees_din <= x"03f84904";
		wait for Clk_period;
		Addr <=  "00110101010010";
		Trees_din <= x"004d358d";
		wait for Clk_period;
		Addr <=  "00110101010011";
		Trees_din <= x"ffad358d";
		wait for Clk_period;
		Addr <=  "00110101010100";
		Trees_din <= x"11046d10";
		wait for Clk_period;
		Addr <=  "00110101010101";
		Trees_din <= x"11043808";
		wait for Clk_period;
		Addr <=  "00110101010110";
		Trees_din <= x"18003b04";
		wait for Clk_period;
		Addr <=  "00110101010111";
		Trees_din <= x"0043358d";
		wait for Clk_period;
		Addr <=  "00110101011000";
		Trees_din <= x"0006358d";
		wait for Clk_period;
		Addr <=  "00110101011001";
		Trees_din <= x"10fad204";
		wait for Clk_period;
		Addr <=  "00110101011010";
		Trees_din <= x"0020358d";
		wait for Clk_period;
		Addr <=  "00110101011011";
		Trees_din <= x"ff83358d";
		wait for Clk_period;
		Addr <=  "00110101011100";
		Trees_din <= x"17000008";
		wait for Clk_period;
		Addr <=  "00110101011101";
		Trees_din <= x"0afc9004";
		wait for Clk_period;
		Addr <=  "00110101011110";
		Trees_din <= x"ffa1358d";
		wait for Clk_period;
		Addr <=  "00110101011111";
		Trees_din <= x"0025358d";
		wait for Clk_period;
		Addr <=  "00110101100000";
		Trees_din <= x"1c003f04";
		wait for Clk_period;
		Addr <=  "00110101100001";
		Trees_din <= x"0071358d";
		wait for Clk_period;
		Addr <=  "00110101100010";
		Trees_din <= x"ffef358d";
		wait for Clk_period;
		Addr <=  "00110101100011";
		Trees_din <= x"000fd330";
		wait for Clk_period;
		Addr <=  "00110101100100";
		Trees_din <= x"0b062528";
		wait for Clk_period;
		Addr <=  "00110101100101";
		Trees_din <= x"0b05671c";
		wait for Clk_period;
		Addr <=  "00110101100110";
		Trees_din <= x"09005d10";
		wait for Clk_period;
		Addr <=  "00110101100111";
		Trees_din <= x"020c6008";
		wait for Clk_period;
		Addr <=  "00110101101000";
		Trees_din <= x"010e6604";
		wait for Clk_period;
		Addr <=  "00110101101001";
		Trees_din <= x"00013699";
		wait for Clk_period;
		Addr <=  "00110101101010";
		Trees_din <= x"ffde3699";
		wait for Clk_period;
		Addr <=  "00110101101011";
		Trees_din <= x"03f8e604";
		wait for Clk_period;
		Addr <=  "00110101101100";
		Trees_din <= x"ffec3699";
		wait for Clk_period;
		Addr <=  "00110101101101";
		Trees_din <= x"ff843699";
		wait for Clk_period;
		Addr <=  "00110101101110";
		Trees_din <= x"0f002404";
		wait for Clk_period;
		Addr <=  "00110101101111";
		Trees_din <= x"ffed3699";
		wait for Clk_period;
		Addr <=  "00110101110000";
		Trees_din <= x"18004604";
		wait for Clk_period;
		Addr <=  "00110101110001";
		Trees_din <= x"00753699";
		wait for Clk_period;
		Addr <=  "00110101110010";
		Trees_din <= x"001e3699";
		wait for Clk_period;
		Addr <=  "00110101110011";
		Trees_din <= x"09005808";
		wait for Clk_period;
		Addr <=  "00110101110100";
		Trees_din <= x"0007fa04";
		wait for Clk_period;
		Addr <=  "00110101110101";
		Trees_din <= x"ffe03699";
		wait for Clk_period;
		Addr <=  "00110101110110";
		Trees_din <= x"00833699";
		wait for Clk_period;
		Addr <=  "00110101110111";
		Trees_din <= x"ffd13699";
		wait for Clk_period;
		Addr <=  "00110101111000";
		Trees_din <= x"12fe3504";
		wait for Clk_period;
		Addr <=  "00110101111001";
		Trees_din <= x"ff853699";
		wait for Clk_period;
		Addr <=  "00110101111010";
		Trees_din <= x"00213699";
		wait for Clk_period;
		Addr <=  "00110101111011";
		Trees_din <= x"0c01bf34";
		wait for Clk_period;
		Addr <=  "00110101111100";
		Trees_din <= x"03f7f020";
		wait for Clk_period;
		Addr <=  "00110101111101";
		Trees_din <= x"0d004710";
		wait for Clk_period;
		Addr <=  "00110101111110";
		Trees_din <= x"13fa3508";
		wait for Clk_period;
		Addr <=  "00110101111111";
		Trees_din <= x"0d000004";
		wait for Clk_period;
		Addr <=  "00110110000000";
		Trees_din <= x"ffe23699";
		wait for Clk_period;
		Addr <=  "00110110000001";
		Trees_din <= x"00613699";
		wait for Clk_period;
		Addr <=  "00110110000010";
		Trees_din <= x"03f63504";
		wait for Clk_period;
		Addr <=  "00110110000011";
		Trees_din <= x"fffa3699";
		wait for Clk_period;
		Addr <=  "00110110000100";
		Trees_din <= x"ff683699";
		wait for Clk_period;
		Addr <=  "00110110000101";
		Trees_din <= x"16037f08";
		wait for Clk_period;
		Addr <=  "00110110000110";
		Trees_din <= x"03f28904";
		wait for Clk_period;
		Addr <=  "00110110000111";
		Trees_din <= x"fff53699";
		wait for Clk_period;
		Addr <=  "00110110001000";
		Trees_din <= x"00823699";
		wait for Clk_period;
		Addr <=  "00110110001001";
		Trees_din <= x"010d4f04";
		wait for Clk_period;
		Addr <=  "00110110001010";
		Trees_din <= x"00443699";
		wait for Clk_period;
		Addr <=  "00110110001011";
		Trees_din <= x"ffed3699";
		wait for Clk_period;
		Addr <=  "00110110001100";
		Trees_din <= x"0105bc0c";
		wait for Clk_period;
		Addr <=  "00110110001101";
		Trees_din <= x"14025804";
		wait for Clk_period;
		Addr <=  "00110110001110";
		Trees_din <= x"006d3699";
		wait for Clk_period;
		Addr <=  "00110110001111";
		Trees_din <= x"16010304";
		wait for Clk_period;
		Addr <=  "00110110010000";
		Trees_din <= x"00133699";
		wait for Clk_period;
		Addr <=  "00110110010001";
		Trees_din <= x"ff8e3699";
		wait for Clk_period;
		Addr <=  "00110110010010";
		Trees_din <= x"08024504";
		wait for Clk_period;
		Addr <=  "00110110010011";
		Trees_din <= x"00893699";
		wait for Clk_period;
		Addr <=  "00110110010100";
		Trees_din <= x"001c3699";
		wait for Clk_period;
		Addr <=  "00110110010101";
		Trees_din <= x"0bf9560c";
		wait for Clk_period;
		Addr <=  "00110110010110";
		Trees_din <= x"1900a808";
		wait for Clk_period;
		Addr <=  "00110110010111";
		Trees_din <= x"1a00af04";
		wait for Clk_period;
		Addr <=  "00110110011000";
		Trees_din <= x"00103699";
		wait for Clk_period;
		Addr <=  "00110110011001";
		Trees_din <= x"00873699";
		wait for Clk_period;
		Addr <=  "00110110011010";
		Trees_din <= x"ffd73699";
		wait for Clk_period;
		Addr <=  "00110110011011";
		Trees_din <= x"0d006b08";
		wait for Clk_period;
		Addr <=  "00110110011100";
		Trees_din <= x"03f5cb04";
		wait for Clk_period;
		Addr <=  "00110110011101";
		Trees_din <= x"ffeb3699";
		wait for Clk_period;
		Addr <=  "00110110011110";
		Trees_din <= x"007e3699";
		wait for Clk_period;
		Addr <=  "00110110011111";
		Trees_din <= x"05f81708";
		wait for Clk_period;
		Addr <=  "00110110100000";
		Trees_din <= x"1500a404";
		wait for Clk_period;
		Addr <=  "00110110100001";
		Trees_din <= x"00493699";
		wait for Clk_period;
		Addr <=  "00110110100010";
		Trees_din <= x"ffdf3699";
		wait for Clk_period;
		Addr <=  "00110110100011";
		Trees_din <= x"18003904";
		wait for Clk_period;
		Addr <=  "00110110100100";
		Trees_din <= x"00363699";
		wait for Clk_period;
		Addr <=  "00110110100101";
		Trees_din <= x"ffd13699";
		wait for Clk_period;
		Addr <=  "00110110100110";
		Trees_din <= x"01164278";
		wait for Clk_period;
		Addr <=  "00110110100111";
		Trees_din <= x"000fd33c";
		wait for Clk_period;
		Addr <=  "00110110101000";
		Trees_din <= x"19008720";
		wait for Clk_period;
		Addr <=  "00110110101001";
		Trees_din <= x"05fb8410";
		wait for Clk_period;
		Addr <=  "00110110101010";
		Trees_din <= x"08001708";
		wait for Clk_period;
		Addr <=  "00110110101011";
		Trees_din <= x"0afced04";
		wait for Clk_period;
		Addr <=  "00110110101100";
		Trees_din <= x"ffad3795";
		wait for Clk_period;
		Addr <=  "00110110101101";
		Trees_din <= x"00603795";
		wait for Clk_period;
		Addr <=  "00110110101110";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00110110101111";
		Trees_din <= x"00273795";
		wait for Clk_period;
		Addr <=  "00110110110000";
		Trees_din <= x"ff7c3795";
		wait for Clk_period;
		Addr <=  "00110110110001";
		Trees_din <= x"0107ac08";
		wait for Clk_period;
		Addr <=  "00110110110010";
		Trees_din <= x"15009404";
		wait for Clk_period;
		Addr <=  "00110110110011";
		Trees_din <= x"ffd63795";
		wait for Clk_period;
		Addr <=  "00110110110100";
		Trees_din <= x"00543795";
		wait for Clk_period;
		Addr <=  "00110110110101";
		Trees_din <= x"0b028704";
		wait for Clk_period;
		Addr <=  "00110110110110";
		Trees_din <= x"00643795";
		wait for Clk_period;
		Addr <=  "00110110110111";
		Trees_din <= x"00013795";
		wait for Clk_period;
		Addr <=  "00110110111000";
		Trees_din <= x"1e007610";
		wait for Clk_period;
		Addr <=  "00110110111001";
		Trees_din <= x"18004808";
		wait for Clk_period;
		Addr <=  "00110110111010";
		Trees_din <= x"18004704";
		wait for Clk_period;
		Addr <=  "00110110111011";
		Trees_din <= x"fffb3795";
		wait for Clk_period;
		Addr <=  "00110110111100";
		Trees_din <= x"00513795";
		wait for Clk_period;
		Addr <=  "00110110111101";
		Trees_din <= x"02005904";
		wait for Clk_period;
		Addr <=  "00110110111110";
		Trees_din <= x"000c3795";
		wait for Clk_period;
		Addr <=  "00110110111111";
		Trees_din <= x"ff8c3795";
		wait for Clk_period;
		Addr <=  "00110111000000";
		Trees_din <= x"1403c908";
		wait for Clk_period;
		Addr <=  "00110111000001";
		Trees_din <= x"02023e04";
		wait for Clk_period;
		Addr <=  "00110111000010";
		Trees_din <= x"ffe93795";
		wait for Clk_period;
		Addr <=  "00110111000011";
		Trees_din <= x"00703795";
		wait for Clk_period;
		Addr <=  "00110111000100";
		Trees_din <= x"ffa93795";
		wait for Clk_period;
		Addr <=  "00110111000101";
		Trees_din <= x"09005a20";
		wait for Clk_period;
		Addr <=  "00110111000110";
		Trees_din <= x"0afb0110";
		wait for Clk_period;
		Addr <=  "00110111000111";
		Trees_din <= x"1a00c508";
		wait for Clk_period;
		Addr <=  "00110111001000";
		Trees_din <= x"0d032504";
		wait for Clk_period;
		Addr <=  "00110111001001";
		Trees_din <= x"00593795";
		wait for Clk_period;
		Addr <=  "00110111001010";
		Trees_din <= x"ffe83795";
		wait for Clk_period;
		Addr <=  "00110111001011";
		Trees_din <= x"1c003104";
		wait for Clk_period;
		Addr <=  "00110111001100";
		Trees_din <= x"000d3795";
		wait for Clk_period;
		Addr <=  "00110111001101";
		Trees_din <= x"ff9b3795";
		wait for Clk_period;
		Addr <=  "00110111001110";
		Trees_din <= x"0c039b08";
		wait for Clk_period;
		Addr <=  "00110111001111";
		Trees_din <= x"0202f304";
		wait for Clk_period;
		Addr <=  "00110111010000";
		Trees_din <= x"00503795";
		wait for Clk_period;
		Addr <=  "00110111010001";
		Trees_din <= x"00183795";
		wait for Clk_period;
		Addr <=  "00110111010010";
		Trees_din <= x"1a00bd04";
		wait for Clk_period;
		Addr <=  "00110111010011";
		Trees_din <= x"00403795";
		wait for Clk_period;
		Addr <=  "00110111010100";
		Trees_din <= x"ffb53795";
		wait for Clk_period;
		Addr <=  "00110111010101";
		Trees_din <= x"1102840c";
		wait for Clk_period;
		Addr <=  "00110111010110";
		Trees_din <= x"1200ea08";
		wait for Clk_period;
		Addr <=  "00110111010111";
		Trees_din <= x"0107ac04";
		wait for Clk_period;
		Addr <=  "00110111011000";
		Trees_din <= x"00333795";
		wait for Clk_period;
		Addr <=  "00110111011001";
		Trees_din <= x"ffb43795";
		wait for Clk_period;
		Addr <=  "00110111011010";
		Trees_din <= x"00613795";
		wait for Clk_period;
		Addr <=  "00110111011011";
		Trees_din <= x"0bfae008";
		wait for Clk_period;
		Addr <=  "00110111011100";
		Trees_din <= x"08014504";
		wait for Clk_period;
		Addr <=  "00110111011101";
		Trees_din <= x"ffd43795";
		wait for Clk_period;
		Addr <=  "00110111011110";
		Trees_din <= x"ff7d3795";
		wait for Clk_period;
		Addr <=  "00110111011111";
		Trees_din <= x"06f4b504";
		wait for Clk_period;
		Addr <=  "00110111100000";
		Trees_din <= x"ffc73795";
		wait for Clk_period;
		Addr <=  "00110111100001";
		Trees_din <= x"001f3795";
		wait for Clk_period;
		Addr <=  "00110111100010";
		Trees_din <= x"09005704";
		wait for Clk_period;
		Addr <=  "00110111100011";
		Trees_din <= x"ffa43795";
		wait for Clk_period;
		Addr <=  "00110111100100";
		Trees_din <= x"fffa3795";
		wait for Clk_period;
		Addr <=  "00110111100101";
		Trees_din <= x"06f34c2c";
		wait for Clk_period;
		Addr <=  "00110111100110";
		Trees_din <= x"0006810c";
		wait for Clk_period;
		Addr <=  "00110111100111";
		Trees_din <= x"0304d308";
		wait for Clk_period;
		Addr <=  "00110111101000";
		Trees_din <= x"05fbbb04";
		wait for Clk_period;
		Addr <=  "00110111101001";
		Trees_din <= x"ff893891";
		wait for Clk_period;
		Addr <=  "00110111101010";
		Trees_din <= x"ffe13891";
		wait for Clk_period;
		Addr <=  "00110111101011";
		Trees_din <= x"002d3891";
		wait for Clk_period;
		Addr <=  "00110111101100";
		Trees_din <= x"03feb01c";
		wait for Clk_period;
		Addr <=  "00110111101101";
		Trees_din <= x"0c02c110";
		wait for Clk_period;
		Addr <=  "00110111101110";
		Trees_din <= x"0c00d708";
		wait for Clk_period;
		Addr <=  "00110111101111";
		Trees_din <= x"09005904";
		wait for Clk_period;
		Addr <=  "00110111110000";
		Trees_din <= x"00513891";
		wait for Clk_period;
		Addr <=  "00110111110001";
		Trees_din <= x"ffd23891";
		wait for Clk_period;
		Addr <=  "00110111110010";
		Trees_din <= x"0203bd04";
		wait for Clk_period;
		Addr <=  "00110111110011";
		Trees_din <= x"00373891";
		wait for Clk_period;
		Addr <=  "00110111110100";
		Trees_din <= x"ffc83891";
		wait for Clk_period;
		Addr <=  "00110111110101";
		Trees_din <= x"01128f08";
		wait for Clk_period;
		Addr <=  "00110111110110";
		Trees_din <= x"1d004004";
		wait for Clk_period;
		Addr <=  "00110111110111";
		Trees_din <= x"000c3891";
		wait for Clk_period;
		Addr <=  "00110111111000";
		Trees_din <= x"007e3891";
		wait for Clk_period;
		Addr <=  "00110111111001";
		Trees_din <= x"ffca3891";
		wait for Clk_period;
		Addr <=  "00110111111010";
		Trees_din <= x"00893891";
		wait for Clk_period;
		Addr <=  "00110111111011";
		Trees_din <= x"0209442c";
		wait for Clk_period;
		Addr <=  "00110111111100";
		Trees_din <= x"02089520";
		wait for Clk_period;
		Addr <=  "00110111111101";
		Trees_din <= x"09005810";
		wait for Clk_period;
		Addr <=  "00110111111110";
		Trees_din <= x"10fb1d08";
		wait for Clk_period;
		Addr <=  "00110111111111";
		Trees_din <= x"10faf104";
		wait for Clk_period;
		Addr <=  "00111000000000";
		Trees_din <= x"00033891";
		wait for Clk_period;
		Addr <=  "00111000000001";
		Trees_din <= x"005a3891";
		wait for Clk_period;
		Addr <=  "00111000000010";
		Trees_din <= x"01019804";
		wait for Clk_period;
		Addr <=  "00111000000011";
		Trees_din <= x"00173891";
		wait for Clk_period;
		Addr <=  "00111000000100";
		Trees_din <= x"ffe73891";
		wait for Clk_period;
		Addr <=  "00111000000101";
		Trees_din <= x"13fef608";
		wait for Clk_period;
		Addr <=  "00111000000110";
		Trees_din <= x"0d000e04";
		wait for Clk_period;
		Addr <=  "00111000000111";
		Trees_din <= x"ffce3891";
		wait for Clk_period;
		Addr <=  "00111000001000";
		Trees_din <= x"00473891";
		wait for Clk_period;
		Addr <=  "00111000001001";
		Trees_din <= x"08018604";
		wait for Clk_period;
		Addr <=  "00111000001010";
		Trees_din <= x"ffdd3891";
		wait for Clk_period;
		Addr <=  "00111000001011";
		Trees_din <= x"00273891";
		wait for Clk_period;
		Addr <=  "00111000001100";
		Trees_din <= x"0b040408";
		wait for Clk_period;
		Addr <=  "00111000001101";
		Trees_din <= x"06f6f704";
		wait for Clk_period;
		Addr <=  "00111000001110";
		Trees_din <= x"00863891";
		wait for Clk_period;
		Addr <=  "00111000001111";
		Trees_din <= x"00183891";
		wait for Clk_period;
		Addr <=  "00111000010000";
		Trees_din <= x"ffd13891";
		wait for Clk_period;
		Addr <=  "00111000010001";
		Trees_din <= x"0c026320";
		wait for Clk_period;
		Addr <=  "00111000010010";
		Trees_din <= x"18004310";
		wait for Clk_period;
		Addr <=  "00111000010011";
		Trees_din <= x"08013908";
		wait for Clk_period;
		Addr <=  "00111000010100";
		Trees_din <= x"0efff404";
		wait for Clk_period;
		Addr <=  "00111000010101";
		Trees_din <= x"ffe63891";
		wait for Clk_period;
		Addr <=  "00111000010110";
		Trees_din <= x"00753891";
		wait for Clk_period;
		Addr <=  "00111000010111";
		Trees_din <= x"1603d304";
		wait for Clk_period;
		Addr <=  "00111000011000";
		Trees_din <= x"ffb93891";
		wait for Clk_period;
		Addr <=  "00111000011001";
		Trees_din <= x"003b3891";
		wait for Clk_period;
		Addr <=  "00111000011010";
		Trees_din <= x"0c00f908";
		wait for Clk_period;
		Addr <=  "00111000011011";
		Trees_din <= x"000fd304";
		wait for Clk_period;
		Addr <=  "00111000011100";
		Trees_din <= x"ff803891";
		wait for Clk_period;
		Addr <=  "00111000011101";
		Trees_din <= x"ffdb3891";
		wait for Clk_period;
		Addr <=  "00111000011110";
		Trees_din <= x"0c01b504";
		wait for Clk_period;
		Addr <=  "00111000011111";
		Trees_din <= x"00453891";
		wait for Clk_period;
		Addr <=  "00111000100000";
		Trees_din <= x"ffc13891";
		wait for Clk_period;
		Addr <=  "00111000100001";
		Trees_din <= x"11031504";
		wait for Clk_period;
		Addr <=  "00111000100010";
		Trees_din <= x"ff7d3891";
		wait for Clk_period;
		Addr <=  "00111000100011";
		Trees_din <= x"fff93891";
		wait for Clk_period;
		Addr <=  "00111000100100";
		Trees_din <= x"000b1e3c";
		wait for Clk_period;
		Addr <=  "00111000100101";
		Trees_din <= x"21000030";
		wait for Clk_period;
		Addr <=  "00111000100110";
		Trees_din <= x"05fe5c18";
		wait for Clk_period;
		Addr <=  "00111000100111";
		Trees_din <= x"020abe10";
		wait for Clk_period;
		Addr <=  "00111000101000";
		Trees_din <= x"010ea208";
		wait for Clk_period;
		Addr <=  "00111000101001";
		Trees_din <= x"19009904";
		wait for Clk_period;
		Addr <=  "00111000101010";
		Trees_din <= x"fff739a5";
		wait for Clk_period;
		Addr <=  "00111000101011";
		Trees_din <= x"002639a5";
		wait for Clk_period;
		Addr <=  "00111000101100";
		Trees_din <= x"12028704";
		wait for Clk_period;
		Addr <=  "00111000101101";
		Trees_din <= x"ff9d39a5";
		wait for Clk_period;
		Addr <=  "00111000101110";
		Trees_din <= x"001639a5";
		wait for Clk_period;
		Addr <=  "00111000101111";
		Trees_din <= x"1900a604";
		wait for Clk_period;
		Addr <=  "00111000110000";
		Trees_din <= x"ff8b39a5";
		wait for Clk_period;
		Addr <=  "00111000110001";
		Trees_din <= x"001439a5";
		wait for Clk_period;
		Addr <=  "00111000110010";
		Trees_din <= x"19009b10";
		wait for Clk_period;
		Addr <=  "00111000110011";
		Trees_din <= x"18004608";
		wait for Clk_period;
		Addr <=  "00111000110100";
		Trees_din <= x"15009904";
		wait for Clk_period;
		Addr <=  "00111000110101";
		Trees_din <= x"005a39a5";
		wait for Clk_period;
		Addr <=  "00111000110110";
		Trees_din <= x"ffcb39a5";
		wait for Clk_period;
		Addr <=  "00111000110111";
		Trees_din <= x"01fcd904";
		wait for Clk_period;
		Addr <=  "00111000111000";
		Trees_din <= x"001539a5";
		wait for Clk_period;
		Addr <=  "00111000111001";
		Trees_din <= x"ff8d39a5";
		wait for Clk_period;
		Addr <=  "00111000111010";
		Trees_din <= x"1d003904";
		wait for Clk_period;
		Addr <=  "00111000111011";
		Trees_din <= x"ffea39a5";
		wait for Clk_period;
		Addr <=  "00111000111100";
		Trees_din <= x"ff8639a5";
		wait for Clk_period;
		Addr <=  "00111000111101";
		Trees_din <= x"01005e04";
		wait for Clk_period;
		Addr <=  "00111000111110";
		Trees_din <= x"003239a5";
		wait for Clk_period;
		Addr <=  "00111000111111";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00111001000000";
		Trees_din <= x"ffde39a5";
		wait for Clk_period;
		Addr <=  "00111001000001";
		Trees_din <= x"ff7c39a5";
		wait for Clk_period;
		Addr <=  "00111001000010";
		Trees_din <= x"18003618";
		wait for Clk_period;
		Addr <=  "00111001000011";
		Trees_din <= x"010db60c";
		wait for Clk_period;
		Addr <=  "00111001000100";
		Trees_din <= x"03f68204";
		wait for Clk_period;
		Addr <=  "00111001000101";
		Trees_din <= x"fff739a5";
		wait for Clk_period;
		Addr <=  "00111001000110";
		Trees_din <= x"000d2304";
		wait for Clk_period;
		Addr <=  "00111001000111";
		Trees_din <= x"001b39a5";
		wait for Clk_period;
		Addr <=  "00111001001000";
		Trees_din <= x"008139a5";
		wait for Clk_period;
		Addr <=  "00111001001001";
		Trees_din <= x"0d00a704";
		wait for Clk_period;
		Addr <=  "00111001001010";
		Trees_din <= x"005139a5";
		wait for Clk_period;
		Addr <=  "00111001001011";
		Trees_din <= x"00100404";
		wait for Clk_period;
		Addr <=  "00111001001100";
		Trees_din <= x"ffa239a5";
		wait for Clk_period;
		Addr <=  "00111001001101";
		Trees_din <= x"000939a5";
		wait for Clk_period;
		Addr <=  "00111001001110";
		Trees_din <= x"1b003618";
		wait for Clk_period;
		Addr <=  "00111001001111";
		Trees_din <= x"1c002a08";
		wait for Clk_period;
		Addr <=  "00111001010000";
		Trees_din <= x"0202b804";
		wait for Clk_period;
		Addr <=  "00111001010001";
		Trees_din <= x"fff539a5";
		wait for Clk_period;
		Addr <=  "00111001010010";
		Trees_din <= x"ff8e39a5";
		wait for Clk_period;
		Addr <=  "00111001010011";
		Trees_din <= x"010f3708";
		wait for Clk_period;
		Addr <=  "00111001010100";
		Trees_din <= x"03fd6504";
		wait for Clk_period;
		Addr <=  "00111001010101";
		Trees_din <= x"ffda39a5";
		wait for Clk_period;
		Addr <=  "00111001010110";
		Trees_din <= x"005a39a5";
		wait for Clk_period;
		Addr <=  "00111001010111";
		Trees_din <= x"0f01a804";
		wait for Clk_period;
		Addr <=  "00111001011000";
		Trees_din <= x"ffde39a5";
		wait for Clk_period;
		Addr <=  "00111001011001";
		Trees_din <= x"005d39a5";
		wait for Clk_period;
		Addr <=  "00111001011010";
		Trees_din <= x"1a00cb10";
		wait for Clk_period;
		Addr <=  "00111001011011";
		Trees_din <= x"0d036508";
		wait for Clk_period;
		Addr <=  "00111001011100";
		Trees_din <= x"11ff1104";
		wait for Clk_period;
		Addr <=  "00111001011101";
		Trees_din <= x"003139a5";
		wait for Clk_period;
		Addr <=  "00111001011110";
		Trees_din <= x"ffed39a5";
		wait for Clk_period;
		Addr <=  "00111001011111";
		Trees_din <= x"09005404";
		wait for Clk_period;
		Addr <=  "00111001100000";
		Trees_din <= x"fff539a5";
		wait for Clk_period;
		Addr <=  "00111001100001";
		Trees_din <= x"004d39a5";
		wait for Clk_period;
		Addr <=  "00111001100010";
		Trees_din <= x"1d004808";
		wait for Clk_period;
		Addr <=  "00111001100011";
		Trees_din <= x"1500ac04";
		wait for Clk_period;
		Addr <=  "00111001100100";
		Trees_din <= x"007139a5";
		wait for Clk_period;
		Addr <=  "00111001100101";
		Trees_din <= x"ffe739a5";
		wait for Clk_period;
		Addr <=  "00111001100110";
		Trees_din <= x"17000204";
		wait for Clk_period;
		Addr <=  "00111001100111";
		Trees_din <= x"ffa239a5";
		wait for Clk_period;
		Addr <=  "00111001101000";
		Trees_din <= x"000f39a5";
		wait for Clk_period;
		Addr <=  "00111001101001";
		Trees_din <= x"000fd32c";
		wait for Clk_period;
		Addr <=  "00111001101010";
		Trees_din <= x"09005d24";
		wait for Clk_period;
		Addr <=  "00111001101011";
		Trees_din <= x"0b06251c";
		wait for Clk_period;
		Addr <=  "00111001101100";
		Trees_din <= x"0b056710";
		wait for Clk_period;
		Addr <=  "00111001101101";
		Trees_din <= x"03fe5108";
		wait for Clk_period;
		Addr <=  "00111001101110";
		Trees_din <= x"0f006804";
		wait for Clk_period;
		Addr <=  "00111001101111";
		Trees_din <= x"ffd43a89";
		wait for Clk_period;
		Addr <=  "00111001110000";
		Trees_din <= x"fffd3a89";
		wait for Clk_period;
		Addr <=  "00111001110001";
		Trees_din <= x"000b5604";
		wait for Clk_period;
		Addr <=  "00111001110010";
		Trees_din <= x"fffe3a89";
		wait for Clk_period;
		Addr <=  "00111001110011";
		Trees_din <= x"00533a89";
		wait for Clk_period;
		Addr <=  "00111001110100";
		Trees_din <= x"12ff0204";
		wait for Clk_period;
		Addr <=  "00111001110101";
		Trees_din <= x"ffdf3a89";
		wait for Clk_period;
		Addr <=  "00111001110110";
		Trees_din <= x"02013704";
		wait for Clk_period;
		Addr <=  "00111001110111";
		Trees_din <= x"ffef3a89";
		wait for Clk_period;
		Addr <=  "00111001111000";
		Trees_din <= x"007a3a89";
		wait for Clk_period;
		Addr <=  "00111001111001";
		Trees_din <= x"06f7d504";
		wait for Clk_period;
		Addr <=  "00111001111010";
		Trees_din <= x"ff973a89";
		wait for Clk_period;
		Addr <=  "00111001111011";
		Trees_din <= x"fffb3a89";
		wait for Clk_period;
		Addr <=  "00111001111100";
		Trees_din <= x"0f002404";
		wait for Clk_period;
		Addr <=  "00111001111101";
		Trees_din <= x"ffed3a89";
		wait for Clk_period;
		Addr <=  "00111001111110";
		Trees_din <= x"00573a89";
		wait for Clk_period;
		Addr <=  "00111001111111";
		Trees_din <= x"09005a34";
		wait for Clk_period;
		Addr <=  "00111010000000";
		Trees_din <= x"11ff5414";
		wait for Clk_period;
		Addr <=  "00111010000001";
		Trees_din <= x"07005308";
		wait for Clk_period;
		Addr <=  "00111010000010";
		Trees_din <= x"0c010a04";
		wait for Clk_period;
		Addr <=  "00111010000011";
		Trees_din <= x"ffb83a89";
		wait for Clk_period;
		Addr <=  "00111010000100";
		Trees_din <= x"00273a89";
		wait for Clk_period;
		Addr <=  "00111010000101";
		Trees_din <= x"00105d04";
		wait for Clk_period;
		Addr <=  "00111010000110";
		Trees_din <= x"fff43a89";
		wait for Clk_period;
		Addr <=  "00111010000111";
		Trees_din <= x"18003b04";
		wait for Clk_period;
		Addr <=  "00111010001000";
		Trees_din <= x"00113a89";
		wait for Clk_period;
		Addr <=  "00111010001001";
		Trees_din <= x"00853a89";
		wait for Clk_period;
		Addr <=  "00111010001010";
		Trees_din <= x"1100c210";
		wait for Clk_period;
		Addr <=  "00111010001011";
		Trees_din <= x"010d4f08";
		wait for Clk_period;
		Addr <=  "00111010001100";
		Trees_din <= x"1004bf04";
		wait for Clk_period;
		Addr <=  "00111010001101";
		Trees_din <= x"00693a89";
		wait for Clk_period;
		Addr <=  "00111010001110";
		Trees_din <= x"ffc13a89";
		wait for Clk_period;
		Addr <=  "00111010001111";
		Trees_din <= x"05f92804";
		wait for Clk_period;
		Addr <=  "00111010010000";
		Trees_din <= x"ffee3a89";
		wait for Clk_period;
		Addr <=  "00111010010001";
		Trees_din <= x"ff8a3a89";
		wait for Clk_period;
		Addr <=  "00111010010010";
		Trees_din <= x"0b046c08";
		wait for Clk_period;
		Addr <=  "00111010010011";
		Trees_din <= x"1403e404";
		wait for Clk_period;
		Addr <=  "00111010010100";
		Trees_din <= x"00253a89";
		wait for Clk_period;
		Addr <=  "00111010010101";
		Trees_din <= x"ffd63a89";
		wait for Clk_period;
		Addr <=  "00111010010110";
		Trees_din <= x"0011cf04";
		wait for Clk_period;
		Addr <=  "00111010010111";
		Trees_din <= x"ffab3a89";
		wait for Clk_period;
		Addr <=  "00111010011000";
		Trees_din <= x"000f3a89";
		wait for Clk_period;
		Addr <=  "00111010011001";
		Trees_din <= x"0bf96e04";
		wait for Clk_period;
		Addr <=  "00111010011010";
		Trees_din <= x"003d3a89";
		wait for Clk_period;
		Addr <=  "00111010011011";
		Trees_din <= x"0b048f0c";
		wait for Clk_period;
		Addr <=  "00111010011100";
		Trees_din <= x"0d010104";
		wait for Clk_period;
		Addr <=  "00111010011101";
		Trees_din <= x"001c3a89";
		wait for Clk_period;
		Addr <=  "00111010011110";
		Trees_din <= x"0800e004";
		wait for Clk_period;
		Addr <=  "00111010011111";
		Trees_din <= x"ffef3a89";
		wait for Clk_period;
		Addr <=  "00111010100000";
		Trees_din <= x"ff8c3a89";
		wait for Clk_period;
		Addr <=  "00111010100001";
		Trees_din <= x"00233a89";
		wait for Clk_period;
		Addr <=  "00111010100010";
		Trees_din <= x"0003aa20";
		wait for Clk_period;
		Addr <=  "00111010100011";
		Trees_din <= x"1b003d10";
		wait for Clk_period;
		Addr <=  "00111010100100";
		Trees_din <= x"08022f08";
		wait for Clk_period;
		Addr <=  "00111010100101";
		Trees_din <= x"03075d04";
		wait for Clk_period;
		Addr <=  "00111010100110";
		Trees_din <= x"ff8d3b85";
		wait for Clk_period;
		Addr <=  "00111010100111";
		Trees_din <= x"fffd3b85";
		wait for Clk_period;
		Addr <=  "00111010101000";
		Trees_din <= x"0afde304";
		wait for Clk_period;
		Addr <=  "00111010101001";
		Trees_din <= x"003f3b85";
		wait for Clk_period;
		Addr <=  "00111010101010";
		Trees_din <= x"ffae3b85";
		wait for Clk_period;
		Addr <=  "00111010101011";
		Trees_din <= x"0700580c";
		wait for Clk_period;
		Addr <=  "00111010101100";
		Trees_din <= x"0c01fd08";
		wait for Clk_period;
		Addr <=  "00111010101101";
		Trees_din <= x"0c012004";
		wait for Clk_period;
		Addr <=  "00111010101110";
		Trees_din <= x"fff03b85";
		wait for Clk_period;
		Addr <=  "00111010101111";
		Trees_din <= x"005e3b85";
		wait for Clk_period;
		Addr <=  "00111010110000";
		Trees_din <= x"ffe63b85";
		wait for Clk_period;
		Addr <=  "00111010110001";
		Trees_din <= x"ffc83b85";
		wait for Clk_period;
		Addr <=  "00111010110010";
		Trees_din <= x"02ffbf24";
		wait for Clk_period;
		Addr <=  "00111010110011";
		Trees_din <= x"06f68b10";
		wait for Clk_period;
		Addr <=  "00111010110100";
		Trees_din <= x"0d03310c";
		wait for Clk_period;
		Addr <=  "00111010110101";
		Trees_din <= x"13f8dd04";
		wait for Clk_period;
		Addr <=  "00111010110110";
		Trees_din <= x"fff03b85";
		wait for Clk_period;
		Addr <=  "00111010110111";
		Trees_din <= x"07005b04";
		wait for Clk_period;
		Addr <=  "00111010111000";
		Trees_din <= x"00753b85";
		wait for Clk_period;
		Addr <=  "00111010111001";
		Trees_din <= x"00103b85";
		wait for Clk_period;
		Addr <=  "00111010111010";
		Trees_din <= x"ffe33b85";
		wait for Clk_period;
		Addr <=  "00111010111011";
		Trees_din <= x"0f003e08";
		wait for Clk_period;
		Addr <=  "00111010111100";
		Trees_din <= x"0b041504";
		wait for Clk_period;
		Addr <=  "00111010111101";
		Trees_din <= x"00663b85";
		wait for Clk_period;
		Addr <=  "00111010111110";
		Trees_din <= x"00013b85";
		wait for Clk_period;
		Addr <=  "00111010111111";
		Trees_din <= x"10f9dc04";
		wait for Clk_period;
		Addr <=  "00111011000000";
		Trees_din <= x"00413b85";
		wait for Clk_period;
		Addr <=  "00111011000001";
		Trees_din <= x"10028704";
		wait for Clk_period;
		Addr <=  "00111011000010";
		Trees_din <= x"ffba3b85";
		wait for Clk_period;
		Addr <=  "00111011000011";
		Trees_din <= x"00173b85";
		wait for Clk_period;
		Addr <=  "00111011000100";
		Trees_din <= x"06f34c1c";
		wait for Clk_period;
		Addr <=  "00111011000101";
		Trees_din <= x"1101fb0c";
		wait for Clk_period;
		Addr <=  "00111011000110";
		Trees_din <= x"0112d608";
		wait for Clk_period;
		Addr <=  "00111011000111";
		Trees_din <= x"1005a904";
		wait for Clk_period;
		Addr <=  "00111011001000";
		Trees_din <= x"005a3b85";
		wait for Clk_period;
		Addr <=  "00111011001001";
		Trees_din <= x"ffd43b85";
		wait for Clk_period;
		Addr <=  "00111011001010";
		Trees_din <= x"ffcd3b85";
		wait for Clk_period;
		Addr <=  "00111011001011";
		Trees_din <= x"0c00cd08";
		wait for Clk_period;
		Addr <=  "00111011001100";
		Trees_din <= x"09005904";
		wait for Clk_period;
		Addr <=  "00111011001101";
		Trees_din <= x"00593b85";
		wait for Clk_period;
		Addr <=  "00111011001110";
		Trees_din <= x"ffd43b85";
		wait for Clk_period;
		Addr <=  "00111011001111";
		Trees_din <= x"0c01df04";
		wait for Clk_period;
		Addr <=  "00111011010000";
		Trees_din <= x"ffaf3b85";
		wait for Clk_period;
		Addr <=  "00111011010001";
		Trees_din <= x"00153b85";
		wait for Clk_period;
		Addr <=  "00111011010010";
		Trees_din <= x"1900a110";
		wait for Clk_period;
		Addr <=  "00111011010011";
		Trees_din <= x"06f3ec08";
		wait for Clk_period;
		Addr <=  "00111011010100";
		Trees_din <= x"10052104";
		wait for Clk_period;
		Addr <=  "00111011010101";
		Trees_din <= x"ffa43b85";
		wait for Clk_period;
		Addr <=  "00111011010110";
		Trees_din <= x"000f3b85";
		wait for Clk_period;
		Addr <=  "00111011010111";
		Trees_din <= x"19009c04";
		wait for Clk_period;
		Addr <=  "00111011011000";
		Trees_din <= x"00043b85";
		wait for Clk_period;
		Addr <=  "00111011011001";
		Trees_din <= x"ffd03b85";
		wait for Clk_period;
		Addr <=  "00111011011010";
		Trees_din <= x"0c033108";
		wait for Clk_period;
		Addr <=  "00111011011011";
		Trees_din <= x"09005004";
		wait for Clk_period;
		Addr <=  "00111011011100";
		Trees_din <= x"fff03b85";
		wait for Clk_period;
		Addr <=  "00111011011101";
		Trees_din <= x"00363b85";
		wait for Clk_period;
		Addr <=  "00111011011110";
		Trees_din <= x"0109bf04";
		wait for Clk_period;
		Addr <=  "00111011011111";
		Trees_din <= x"00203b85";
		wait for Clk_period;
		Addr <=  "00111011100000";
		Trees_din <= x"ff993b85";
		wait for Clk_period;
		Addr <=  "00111011100001";
		Trees_din <= x"000f6f34";
		wait for Clk_period;
		Addr <=  "00111011100010";
		Trees_din <= x"09005d28";
		wait for Clk_period;
		Addr <=  "00111011100011";
		Trees_din <= x"21000020";
		wait for Clk_period;
		Addr <=  "00111011100100";
		Trees_din <= x"15008c10";
		wait for Clk_period;
		Addr <=  "00111011100101";
		Trees_din <= x"0401a508";
		wait for Clk_period;
		Addr <=  "00111011100110";
		Trees_din <= x"0c018304";
		wait for Clk_period;
		Addr <=  "00111011100111";
		Trees_din <= x"ffac3c59";
		wait for Clk_period;
		Addr <=  "00111011101000";
		Trees_din <= x"fff43c59";
		wait for Clk_period;
		Addr <=  "00111011101001";
		Trees_din <= x"00025704";
		wait for Clk_period;
		Addr <=  "00111011101010";
		Trees_din <= x"ffb93c59";
		wait for Clk_period;
		Addr <=  "00111011101011";
		Trees_din <= x"00413c59";
		wait for Clk_period;
		Addr <=  "00111011101100";
		Trees_din <= x"09005808";
		wait for Clk_period;
		Addr <=  "00111011101101";
		Trees_din <= x"0e020504";
		wait for Clk_period;
		Addr <=  "00111011101110";
		Trees_din <= x"ffe83c59";
		wait for Clk_period;
		Addr <=  "00111011101111";
		Trees_din <= x"00163c59";
		wait for Clk_period;
		Addr <=  "00111011110000";
		Trees_din <= x"00054504";
		wait for Clk_period;
		Addr <=  "00111011110001";
		Trees_din <= x"ffa03c59";
		wait for Clk_period;
		Addr <=  "00111011110010";
		Trees_din <= x"00433c59";
		wait for Clk_period;
		Addr <=  "00111011110011";
		Trees_din <= x"04012004";
		wait for Clk_period;
		Addr <=  "00111011110100";
		Trees_din <= x"ffa53c59";
		wait for Clk_period;
		Addr <=  "00111011110101";
		Trees_din <= x"000d3c59";
		wait for Clk_period;
		Addr <=  "00111011110110";
		Trees_din <= x"0f002404";
		wait for Clk_period;
		Addr <=  "00111011110111";
		Trees_din <= x"fff33c59";
		wait for Clk_period;
		Addr <=  "00111011111000";
		Trees_din <= x"0d00ef04";
		wait for Clk_period;
		Addr <=  "00111011111001";
		Trees_din <= x"005f3c59";
		wait for Clk_period;
		Addr <=  "00111011111010";
		Trees_din <= x"00193c59";
		wait for Clk_period;
		Addr <=  "00111011111011";
		Trees_din <= x"04fba420";
		wait for Clk_period;
		Addr <=  "00111011111100";
		Trees_din <= x"0af7a508";
		wait for Clk_period;
		Addr <=  "00111011111101";
		Trees_din <= x"15008704";
		wait for Clk_period;
		Addr <=  "00111011111110";
		Trees_din <= x"fffe3c59";
		wait for Clk_period;
		Addr <=  "00111011111111";
		Trees_din <= x"00703c59";
		wait for Clk_period;
		Addr <=  "00111100000000";
		Trees_din <= x"06fab310";
		wait for Clk_period;
		Addr <=  "00111100000001";
		Trees_din <= x"08000a08";
		wait for Clk_period;
		Addr <=  "00111100000010";
		Trees_din <= x"0afaf604";
		wait for Clk_period;
		Addr <=  "00111100000011";
		Trees_din <= x"fffd3c59";
		wait for Clk_period;
		Addr <=  "00111100000100";
		Trees_din <= x"005e3c59";
		wait for Clk_period;
		Addr <=  "00111100000101";
		Trees_din <= x"03fb9304";
		wait for Clk_period;
		Addr <=  "00111100000110";
		Trees_din <= x"fffc3c59";
		wait for Clk_period;
		Addr <=  "00111100000111";
		Trees_din <= x"ffba3c59";
		wait for Clk_period;
		Addr <=  "00111100001000";
		Trees_din <= x"02ffb904";
		wait for Clk_period;
		Addr <=  "00111100001001";
		Trees_din <= x"ffdd3c59";
		wait for Clk_period;
		Addr <=  "00111100001010";
		Trees_din <= x"006e3c59";
		wait for Clk_period;
		Addr <=  "00111100001011";
		Trees_din <= x"00146010";
		wait for Clk_period;
		Addr <=  "00111100001100";
		Trees_din <= x"0af7ba04";
		wait for Clk_period;
		Addr <=  "00111100001101";
		Trees_din <= x"ffc53c59";
		wait for Clk_period;
		Addr <=  "00111100001110";
		Trees_din <= x"01ff4304";
		wait for Clk_period;
		Addr <=  "00111100001111";
		Trees_din <= x"ffe13c59";
		wait for Clk_period;
		Addr <=  "00111100010000";
		Trees_din <= x"010f7404";
		wait for Clk_period;
		Addr <=  "00111100010001";
		Trees_din <= x"00843c59";
		wait for Clk_period;
		Addr <=  "00111100010010";
		Trees_din <= x"00013c59";
		wait for Clk_period;
		Addr <=  "00111100010011";
		Trees_din <= x"06f68504";
		wait for Clk_period;
		Addr <=  "00111100010100";
		Trees_din <= x"001e3c59";
		wait for Clk_period;
		Addr <=  "00111100010101";
		Trees_din <= x"ffa33c59";
		wait for Clk_period;
		Addr <=  "00111100010110";
		Trees_din <= x"000f6f2c";
		wait for Clk_period;
		Addr <=  "00111100010111";
		Trees_din <= x"03f5ed08";
		wait for Clk_period;
		Addr <=  "00111100011000";
		Trees_din <= x"17000004";
		wait for Clk_period;
		Addr <=  "00111100011001";
		Trees_din <= x"000f3d45";
		wait for Clk_period;
		Addr <=  "00111100011010";
		Trees_din <= x"ff953d45";
		wait for Clk_period;
		Addr <=  "00111100011011";
		Trees_din <= x"09005d18";
		wait for Clk_period;
		Addr <=  "00111100011100";
		Trees_din <= x"16000108";
		wait for Clk_period;
		Addr <=  "00111100011101";
		Trees_din <= x"02004a04";
		wait for Clk_period;
		Addr <=  "00111100011110";
		Trees_din <= x"fff23d45";
		wait for Clk_period;
		Addr <=  "00111100011111";
		Trees_din <= x"ffa53d45";
		wait for Clk_period;
		Addr <=  "00111100100000";
		Trees_din <= x"0d003008";
		wait for Clk_period;
		Addr <=  "00111100100001";
		Trees_din <= x"15008b04";
		wait for Clk_period;
		Addr <=  "00111100100010";
		Trees_din <= x"ffd93d45";
		wait for Clk_period;
		Addr <=  "00111100100011";
		Trees_din <= x"00433d45";
		wait for Clk_period;
		Addr <=  "00111100100100";
		Trees_din <= x"0103e604";
		wait for Clk_period;
		Addr <=  "00111100100101";
		Trees_din <= x"000d3d45";
		wait for Clk_period;
		Addr <=  "00111100100110";
		Trees_din <= x"ffeb3d45";
		wait for Clk_period;
		Addr <=  "00111100100111";
		Trees_din <= x"0f002404";
		wait for Clk_period;
		Addr <=  "00111100101000";
		Trees_din <= x"fff93d45";
		wait for Clk_period;
		Addr <=  "00111100101001";
		Trees_din <= x"0d00ef04";
		wait for Clk_period;
		Addr <=  "00111100101010";
		Trees_din <= x"005c3d45";
		wait for Clk_period;
		Addr <=  "00111100101011";
		Trees_din <= x"00183d45";
		wait for Clk_period;
		Addr <=  "00111100101100";
		Trees_din <= x"1b003828";
		wait for Clk_period;
		Addr <=  "00111100101101";
		Trees_din <= x"06f4800c";
		wait for Clk_period;
		Addr <=  "00111100101110";
		Trees_din <= x"01110604";
		wait for Clk_period;
		Addr <=  "00111100101111";
		Trees_din <= x"007a3d45";
		wait for Clk_period;
		Addr <=  "00111100110000";
		Trees_din <= x"09005404";
		wait for Clk_period;
		Addr <=  "00111100110001";
		Trees_din <= x"ffbe3d45";
		wait for Clk_period;
		Addr <=  "00111100110010";
		Trees_din <= x"00223d45";
		wait for Clk_period;
		Addr <=  "00111100110011";
		Trees_din <= x"18003b10";
		wait for Clk_period;
		Addr <=  "00111100110100";
		Trees_din <= x"0f016808";
		wait for Clk_period;
		Addr <=  "00111100110101";
		Trees_din <= x"010c6804";
		wait for Clk_period;
		Addr <=  "00111100110110";
		Trees_din <= x"002e3d45";
		wait for Clk_period;
		Addr <=  "00111100110111";
		Trees_din <= x"ffc83d45";
		wait for Clk_period;
		Addr <=  "00111100111000";
		Trees_din <= x"04f68004";
		wait for Clk_period;
		Addr <=  "00111100111001";
		Trees_din <= x"00123d45";
		wait for Clk_period;
		Addr <=  "00111100111010";
		Trees_din <= x"00703d45";
		wait for Clk_period;
		Addr <=  "00111100111011";
		Trees_din <= x"0bf95804";
		wait for Clk_period;
		Addr <=  "00111100111100";
		Trees_din <= x"004f3d45";
		wait for Clk_period;
		Addr <=  "00111100111101";
		Trees_din <= x"0bfb0c04";
		wait for Clk_period;
		Addr <=  "00111100111110";
		Trees_din <= x"ff933d45";
		wait for Clk_period;
		Addr <=  "00111100111111";
		Trees_din <= x"ffec3d45";
		wait for Clk_period;
		Addr <=  "00111101000000";
		Trees_din <= x"1e006b0c";
		wait for Clk_period;
		Addr <=  "00111101000001";
		Trees_din <= x"1200b308";
		wait for Clk_period;
		Addr <=  "00111101000010";
		Trees_din <= x"0d02ee04";
		wait for Clk_period;
		Addr <=  "00111101000011";
		Trees_din <= x"004f3d45";
		wait for Clk_period;
		Addr <=  "00111101000100";
		Trees_din <= x"ffd13d45";
		wait for Clk_period;
		Addr <=  "00111101000101";
		Trees_din <= x"00883d45";
		wait for Clk_period;
		Addr <=  "00111101000110";
		Trees_din <= x"11ff1108";
		wait for Clk_period;
		Addr <=  "00111101000111";
		Trees_din <= x"03f2f604";
		wait for Clk_period;
		Addr <=  "00111101001000";
		Trees_din <= x"ffe33d45";
		wait for Clk_period;
		Addr <=  "00111101001001";
		Trees_din <= x"00693d45";
		wait for Clk_period;
		Addr <=  "00111101001010";
		Trees_din <= x"06f57f08";
		wait for Clk_period;
		Addr <=  "00111101001011";
		Trees_din <= x"05fc0a04";
		wait for Clk_period;
		Addr <=  "00111101001100";
		Trees_din <= x"ffd23d45";
		wait for Clk_period;
		Addr <=  "00111101001101";
		Trees_din <= x"002f3d45";
		wait for Clk_period;
		Addr <=  "00111101001110";
		Trees_din <= x"07005b04";
		wait for Clk_period;
		Addr <=  "00111101001111";
		Trees_din <= x"003a3d45";
		wait for Clk_period;
		Addr <=  "00111101010000";
		Trees_din <= x"ffd73d45";
		wait for Clk_period;
		Addr <=  "00111101010001";
		Trees_din <= x"00079050";
		wait for Clk_period;
		Addr <=  "00111101010010";
		Trees_din <= x"03fe251c";
		wait for Clk_period;
		Addr <=  "00111101010011";
		Trees_din <= x"17012b0c";
		wait for Clk_period;
		Addr <=  "00111101010100";
		Trees_din <= x"04ff0108";
		wait for Clk_period;
		Addr <=  "00111101010101";
		Trees_din <= x"16009f04";
		wait for Clk_period;
		Addr <=  "00111101010110";
		Trees_din <= x"00203e81";
		wait for Clk_period;
		Addr <=  "00111101010111";
		Trees_din <= x"ffb03e81";
		wait for Clk_period;
		Addr <=  "00111101011000";
		Trees_din <= x"ff8c3e81";
		wait for Clk_period;
		Addr <=  "00111101011001";
		Trees_din <= x"0f000c04";
		wait for Clk_period;
		Addr <=  "00111101011010";
		Trees_din <= x"ffa43e81";
		wait for Clk_period;
		Addr <=  "00111101011011";
		Trees_din <= x"11021508";
		wait for Clk_period;
		Addr <=  "00111101011100";
		Trees_din <= x"08007104";
		wait for Clk_period;
		Addr <=  "00111101011101";
		Trees_din <= x"005f3e81";
		wait for Clk_period;
		Addr <=  "00111101011110";
		Trees_din <= x"ffff3e81";
		wait for Clk_period;
		Addr <=  "00111101011111";
		Trees_din <= x"ffd93e81";
		wait for Clk_period;
		Addr <=  "00111101100000";
		Trees_din <= x"1201f61c";
		wait for Clk_period;
		Addr <=  "00111101100001";
		Trees_din <= x"0e021e10";
		wait for Clk_period;
		Addr <=  "00111101100010";
		Trees_din <= x"16037108";
		wait for Clk_period;
		Addr <=  "00111101100011";
		Trees_din <= x"06f77604";
		wait for Clk_period;
		Addr <=  "00111101100100";
		Trees_din <= x"ff943e81";
		wait for Clk_period;
		Addr <=  "00111101100101";
		Trees_din <= x"ffe83e81";
		wait for Clk_period;
		Addr <=  "00111101100110";
		Trees_din <= x"09005304";
		wait for Clk_period;
		Addr <=  "00111101100111";
		Trees_din <= x"ffc93e81";
		wait for Clk_period;
		Addr <=  "00111101101000";
		Trees_din <= x"002f3e81";
		wait for Clk_period;
		Addr <=  "00111101101001";
		Trees_din <= x"14014e04";
		wait for Clk_period;
		Addr <=  "00111101101010";
		Trees_din <= x"ffd53e81";
		wait for Clk_period;
		Addr <=  "00111101101011";
		Trees_din <= x"1c003404";
		wait for Clk_period;
		Addr <=  "00111101101100";
		Trees_din <= x"00633e81";
		wait for Clk_period;
		Addr <=  "00111101101101";
		Trees_din <= x"00013e81";
		wait for Clk_period;
		Addr <=  "00111101101110";
		Trees_din <= x"1002880c";
		wait for Clk_period;
		Addr <=  "00111101101111";
		Trees_din <= x"07004f04";
		wait for Clk_period;
		Addr <=  "00111101110000";
		Trees_din <= x"00453e81";
		wait for Clk_period;
		Addr <=  "00111101110001";
		Trees_din <= x"05fcbb04";
		wait for Clk_period;
		Addr <=  "00111101110010";
		Trees_din <= x"ffb33e81";
		wait for Clk_period;
		Addr <=  "00111101110011";
		Trees_din <= x"001a3e81";
		wait for Clk_period;
		Addr <=  "00111101110100";
		Trees_din <= x"1b003004";
		wait for Clk_period;
		Addr <=  "00111101110101";
		Trees_din <= x"007b3e81";
		wait for Clk_period;
		Addr <=  "00111101110110";
		Trees_din <= x"15008704";
		wait for Clk_period;
		Addr <=  "00111101110111";
		Trees_din <= x"005a3e81";
		wait for Clk_period;
		Addr <=  "00111101111000";
		Trees_din <= x"ffcf3e81";
		wait for Clk_period;
		Addr <=  "00111101111001";
		Trees_din <= x"04ff5734";
		wait for Clk_period;
		Addr <=  "00111101111010";
		Trees_din <= x"08001514";
		wait for Clk_period;
		Addr <=  "00111101111011";
		Trees_din <= x"06f96f0c";
		wait for Clk_period;
		Addr <=  "00111101111100";
		Trees_din <= x"01139008";
		wait for Clk_period;
		Addr <=  "00111101111101";
		Trees_din <= x"0f003004";
		wait for Clk_period;
		Addr <=  "00111101111110";
		Trees_din <= x"00033e81";
		wait for Clk_period;
		Addr <=  "00111101111111";
		Trees_din <= x"00553e81";
		wait for Clk_period;
		Addr <=  "00111110000000";
		Trees_din <= x"ffcc3e81";
		wait for Clk_period;
		Addr <=  "00111110000001";
		Trees_din <= x"05fa9804";
		wait for Clk_period;
		Addr <=  "00111110000010";
		Trees_din <= x"ff943e81";
		wait for Clk_period;
		Addr <=  "00111110000011";
		Trees_din <= x"00183e81";
		wait for Clk_period;
		Addr <=  "00111110000100";
		Trees_din <= x"06f5c710";
		wait for Clk_period;
		Addr <=  "00111110000101";
		Trees_din <= x"1f000008";
		wait for Clk_period;
		Addr <=  "00111110000110";
		Trees_din <= x"00105d04";
		wait for Clk_period;
		Addr <=  "00111110000111";
		Trees_din <= x"ffce3e81";
		wait for Clk_period;
		Addr <=  "00111110001000";
		Trees_din <= x"00013e81";
		wait for Clk_period;
		Addr <=  "00111110001001";
		Trees_din <= x"11fec504";
		wait for Clk_period;
		Addr <=  "00111110001010";
		Trees_din <= x"ffc73e81";
		wait for Clk_period;
		Addr <=  "00111110001011";
		Trees_din <= x"003f3e81";
		wait for Clk_period;
		Addr <=  "00111110001100";
		Trees_din <= x"06f63b08";
		wait for Clk_period;
		Addr <=  "00111110001101";
		Trees_din <= x"01065e04";
		wait for Clk_period;
		Addr <=  "00111110001110";
		Trees_din <= x"ffe13e81";
		wait for Clk_period;
		Addr <=  "00111110001111";
		Trees_din <= x"00573e81";
		wait for Clk_period;
		Addr <=  "00111110010000";
		Trees_din <= x"0d00ef04";
		wait for Clk_period;
		Addr <=  "00111110010001";
		Trees_din <= x"001b3e81";
		wait for Clk_period;
		Addr <=  "00111110010010";
		Trees_din <= x"fff33e81";
		wait for Clk_period;
		Addr <=  "00111110010011";
		Trees_din <= x"21000018";
		wait for Clk_period;
		Addr <=  "00111110010100";
		Trees_din <= x"10056f10";
		wait for Clk_period;
		Addr <=  "00111110010101";
		Trees_din <= x"18003d08";
		wait for Clk_period;
		Addr <=  "00111110010110";
		Trees_din <= x"18003b04";
		wait for Clk_period;
		Addr <=  "00111110010111";
		Trees_din <= x"002a3e81";
		wait for Clk_period;
		Addr <=  "00111110011000";
		Trees_din <= x"ffab3e81";
		wait for Clk_period;
		Addr <=  "00111110011001";
		Trees_din <= x"1c004d04";
		wait for Clk_period;
		Addr <=  "00111110011010";
		Trees_din <= x"00673e81";
		wait for Clk_period;
		Addr <=  "00111110011011";
		Trees_din <= x"ffcc3e81";
		wait for Clk_period;
		Addr <=  "00111110011100";
		Trees_din <= x"05fc9304";
		wait for Clk_period;
		Addr <=  "00111110011101";
		Trees_din <= x"00023e81";
		wait for Clk_period;
		Addr <=  "00111110011110";
		Trees_din <= x"ffb73e81";
		wait for Clk_period;
		Addr <=  "00111110011111";
		Trees_din <= x"ffc93e81";
		wait for Clk_period;
		Addr <=  "00111110100000";
		Trees_din <= x"0009b148";
		wait for Clk_period;
		Addr <=  "00111110100001";
		Trees_din <= x"16015b1c";
		wait for Clk_period;
		Addr <=  "00111110100010";
		Trees_din <= x"1201ea08";
		wait for Clk_period;
		Addr <=  "00111110100011";
		Trees_din <= x"0afa1a04";
		wait for Clk_period;
		Addr <=  "00111110100100";
		Trees_din <= x"00123fad";
		wait for Clk_period;
		Addr <=  "00111110100101";
		Trees_din <= x"ff813fad";
		wait for Clk_period;
		Addr <=  "00111110100110";
		Trees_din <= x"0007cf0c";
		wait for Clk_period;
		Addr <=  "00111110100111";
		Trees_din <= x"07005504";
		wait for Clk_period;
		Addr <=  "00111110101000";
		Trees_din <= x"ffd13fad";
		wait for Clk_period;
		Addr <=  "00111110101001";
		Trees_din <= x"09005404";
		wait for Clk_period;
		Addr <=  "00111110101010";
		Trees_din <= x"005f3fad";
		wait for Clk_period;
		Addr <=  "00111110101011";
		Trees_din <= x"fff43fad";
		wait for Clk_period;
		Addr <=  "00111110101100";
		Trees_din <= x"09005804";
		wait for Clk_period;
		Addr <=  "00111110101101";
		Trees_din <= x"ff993fad";
		wait for Clk_period;
		Addr <=  "00111110101110";
		Trees_din <= x"fff93fad";
		wait for Clk_period;
		Addr <=  "00111110101111";
		Trees_din <= x"05fe9620";
		wait for Clk_period;
		Addr <=  "00111110110000";
		Trees_din <= x"06f64110";
		wait for Clk_period;
		Addr <=  "00111110110001";
		Trees_din <= x"05fb6b08";
		wait for Clk_period;
		Addr <=  "00111110110010";
		Trees_din <= x"0f00b004";
		wait for Clk_period;
		Addr <=  "00111110110011";
		Trees_din <= x"002a3fad";
		wait for Clk_period;
		Addr <=  "00111110110100";
		Trees_din <= x"ffb33fad";
		wait for Clk_period;
		Addr <=  "00111110110101";
		Trees_din <= x"0d030504";
		wait for Clk_period;
		Addr <=  "00111110110110";
		Trees_din <= x"005c3fad";
		wait for Clk_period;
		Addr <=  "00111110110111";
		Trees_din <= x"ffe33fad";
		wait for Clk_period;
		Addr <=  "00111110111000";
		Trees_din <= x"0f00ab08";
		wait for Clk_period;
		Addr <=  "00111110111001";
		Trees_din <= x"08005a04";
		wait for Clk_period;
		Addr <=  "00111110111010";
		Trees_din <= x"00103fad";
		wait for Clk_period;
		Addr <=  "00111110111011";
		Trees_din <= x"ff9a3fad";
		wait for Clk_period;
		Addr <=  "00111110111100";
		Trees_din <= x"0801ca04";
		wait for Clk_period;
		Addr <=  "00111110111101";
		Trees_din <= x"ffea3fad";
		wait for Clk_period;
		Addr <=  "00111110111110";
		Trees_din <= x"004d3fad";
		wait for Clk_period;
		Addr <=  "00111110111111";
		Trees_din <= x"06fa5b08";
		wait for Clk_period;
		Addr <=  "00111111000000";
		Trees_din <= x"1b003e04";
		wait for Clk_period;
		Addr <=  "00111111000001";
		Trees_din <= x"ff843fad";
		wait for Clk_period;
		Addr <=  "00111111000010";
		Trees_din <= x"fff73fad";
		wait for Clk_period;
		Addr <=  "00111111000011";
		Trees_din <= x"002f3fad";
		wait for Clk_period;
		Addr <=  "00111111000100";
		Trees_din <= x"18003614";
		wait for Clk_period;
		Addr <=  "00111111000101";
		Trees_din <= x"01087504";
		wait for Clk_period;
		Addr <=  "00111111000110";
		Trees_din <= x"006b3fad";
		wait for Clk_period;
		Addr <=  "00111111000111";
		Trees_din <= x"0206700c";
		wait for Clk_period;
		Addr <=  "00111111001000";
		Trees_din <= x"000d2304";
		wait for Clk_period;
		Addr <=  "00111111001001";
		Trees_din <= x"ffda3fad";
		wait for Clk_period;
		Addr <=  "00111111001010";
		Trees_din <= x"10028604";
		wait for Clk_period;
		Addr <=  "00111111001011";
		Trees_din <= x"006b3fad";
		wait for Clk_period;
		Addr <=  "00111111001100";
		Trees_din <= x"00033fad";
		wait for Clk_period;
		Addr <=  "00111111001101";
		Trees_din <= x"ffba3fad";
		wait for Clk_period;
		Addr <=  "00111111001110";
		Trees_din <= x"1e005c20";
		wait for Clk_period;
		Addr <=  "00111111001111";
		Trees_din <= x"10028810";
		wait for Clk_period;
		Addr <=  "00111111010000";
		Trees_din <= x"010e6608";
		wait for Clk_period;
		Addr <=  "00111111010001";
		Trees_din <= x"07005704";
		wait for Clk_period;
		Addr <=  "00111111010010";
		Trees_din <= x"ff9d3fad";
		wait for Clk_period;
		Addr <=  "00111111010011";
		Trees_din <= x"00113fad";
		wait for Clk_period;
		Addr <=  "00111111010100";
		Trees_din <= x"04fad304";
		wait for Clk_period;
		Addr <=  "00111111010101";
		Trees_din <= x"fffd3fad";
		wait for Clk_period;
		Addr <=  "00111111010110";
		Trees_din <= x"00423fad";
		wait for Clk_period;
		Addr <=  "00111111010111";
		Trees_din <= x"1701c508";
		wait for Clk_period;
		Addr <=  "00111111011000";
		Trees_din <= x"010d4f04";
		wait for Clk_period;
		Addr <=  "00111111011001";
		Trees_din <= x"00783fad";
		wait for Clk_period;
		Addr <=  "00111111011010";
		Trees_din <= x"ffee3fad";
		wait for Clk_period;
		Addr <=  "00111111011011";
		Trees_din <= x"1900a104";
		wait for Clk_period;
		Addr <=  "00111111011100";
		Trees_din <= x"ff983fad";
		wait for Clk_period;
		Addr <=  "00111111011101";
		Trees_din <= x"000a3fad";
		wait for Clk_period;
		Addr <=  "00111111011110";
		Trees_din <= x"11046d10";
		wait for Clk_period;
		Addr <=  "00111111011111";
		Trees_din <= x"05fc2208";
		wait for Clk_period;
		Addr <=  "00111111100000";
		Trees_din <= x"0a028604";
		wait for Clk_period;
		Addr <=  "00111111100001";
		Trees_din <= x"fff03fad";
		wait for Clk_period;
		Addr <=  "00111111100010";
		Trees_din <= x"00183fad";
		wait for Clk_period;
		Addr <=  "00111111100011";
		Trees_din <= x"09005704";
		wait for Clk_period;
		Addr <=  "00111111100100";
		Trees_din <= x"00353fad";
		wait for Clk_period;
		Addr <=  "00111111100101";
		Trees_din <= x"fff83fad";
		wait for Clk_period;
		Addr <=  "00111111100110";
		Trees_din <= x"19008804";
		wait for Clk_period;
		Addr <=  "00111111100111";
		Trees_din <= x"ffe63fad";
		wait for Clk_period;
		Addr <=  "00111111101000";
		Trees_din <= x"17000004";
		wait for Clk_period;
		Addr <=  "00111111101001";
		Trees_din <= x"fff93fad";
		wait for Clk_period;
		Addr <=  "00111111101010";
		Trees_din <= x"00703fad";
		wait for Clk_period;
		Addr <=  "00111111101011";
		Trees_din <= x"000bca40";
		wait for Clk_period;
		Addr <=  "00111111101100";
		Trees_din <= x"1f000838";
		wait for Clk_period;
		Addr <=  "00111111101101";
		Trees_din <= x"19008a18";
		wait for Clk_period;
		Addr <=  "00111111101110";
		Trees_din <= x"04ff7608";
		wait for Clk_period;
		Addr <=  "00111111101111";
		Trees_din <= x"01017504";
		wait for Clk_period;
		Addr <=  "00111111110000";
		Trees_din <= x"fff140a9";
		wait for Clk_period;
		Addr <=  "00111111110001";
		Trees_din <= x"ff8640a9";
		wait for Clk_period;
		Addr <=  "00111111110010";
		Trees_din <= x"0e01d208";
		wait for Clk_period;
		Addr <=  "00111111110011";
		Trees_din <= x"1d005504";
		wait for Clk_period;
		Addr <=  "00111111110100";
		Trees_din <= x"ffbd40a9";
		wait for Clk_period;
		Addr <=  "00111111110101";
		Trees_din <= x"003d40a9";
		wait for Clk_period;
		Addr <=  "00111111110110";
		Trees_din <= x"1d005304";
		wait for Clk_period;
		Addr <=  "00111111110111";
		Trees_din <= x"005040a9";
		wait for Clk_period;
		Addr <=  "00111111111000";
		Trees_din <= x"ffec40a9";
		wait for Clk_period;
		Addr <=  "00111111111001";
		Trees_din <= x"18003d10";
		wait for Clk_period;
		Addr <=  "00111111111010";
		Trees_din <= x"0801aa08";
		wait for Clk_period;
		Addr <=  "00111111111011";
		Trees_din <= x"0afb1a04";
		wait for Clk_period;
		Addr <=  "00111111111100";
		Trees_din <= x"000a40a9";
		wait for Clk_period;
		Addr <=  "00111111111101";
		Trees_din <= x"ffa140a9";
		wait for Clk_period;
		Addr <=  "00111111111110";
		Trees_din <= x"0d010d04";
		wait for Clk_period;
		Addr <=  "00111111111111";
		Trees_din <= x"ffbd40a9";
		wait for Clk_period;
		Addr <=  "01000000000000";
		Trees_din <= x"002b40a9";
		wait for Clk_period;
		Addr <=  "01000000000001";
		Trees_din <= x"0005c708";
		wait for Clk_period;
		Addr <=  "01000000000010";
		Trees_din <= x"08022704";
		wait for Clk_period;
		Addr <=  "01000000000011";
		Trees_din <= x"ffdb40a9";
		wait for Clk_period;
		Addr <=  "01000000000100";
		Trees_din <= x"002b40a9";
		wait for Clk_period;
		Addr <=  "01000000000101";
		Trees_din <= x"21000004";
		wait for Clk_period;
		Addr <=  "01000000000110";
		Trees_din <= x"002d40a9";
		wait for Clk_period;
		Addr <=  "01000000000111";
		Trees_din <= x"ffc340a9";
		wait for Clk_period;
		Addr <=  "01000000001000";
		Trees_din <= x"06f4cb04";
		wait for Clk_period;
		Addr <=  "01000000001001";
		Trees_din <= x"fff440a9";
		wait for Clk_period;
		Addr <=  "01000000001010";
		Trees_din <= x"ff9840a9";
		wait for Clk_period;
		Addr <=  "01000000001011";
		Trees_din <= x"03fd6530";
		wait for Clk_period;
		Addr <=  "01000000001100";
		Trees_din <= x"0bf93b10";
		wait for Clk_period;
		Addr <=  "01000000001101";
		Trees_din <= x"1c002904";
		wait for Clk_period;
		Addr <=  "01000000001110";
		Trees_din <= x"ffc540a9";
		wait for Clk_period;
		Addr <=  "01000000001111";
		Trees_din <= x"07005b08";
		wait for Clk_period;
		Addr <=  "01000000010000";
		Trees_din <= x"04f84b04";
		wait for Clk_period;
		Addr <=  "01000000010001";
		Trees_din <= x"000e40a9";
		wait for Clk_period;
		Addr <=  "01000000010010";
		Trees_din <= x"007e40a9";
		wait for Clk_period;
		Addr <=  "01000000010011";
		Trees_din <= x"ffed40a9";
		wait for Clk_period;
		Addr <=  "01000000010100";
		Trees_din <= x"1d004d10";
		wait for Clk_period;
		Addr <=  "01000000010101";
		Trees_din <= x"1d004c08";
		wait for Clk_period;
		Addr <=  "01000000010110";
		Trees_din <= x"18003604";
		wait for Clk_period;
		Addr <=  "01000000010111";
		Trees_din <= x"003540a9";
		wait for Clk_period;
		Addr <=  "01000000011000";
		Trees_din <= x"fff940a9";
		wait for Clk_period;
		Addr <=  "01000000011001";
		Trees_din <= x"0205dc04";
		wait for Clk_period;
		Addr <=  "01000000011010";
		Trees_din <= x"ff8a40a9";
		wait for Clk_period;
		Addr <=  "01000000011011";
		Trees_din <= x"000240a9";
		wait for Clk_period;
		Addr <=  "01000000011100";
		Trees_din <= x"0a024a08";
		wait for Clk_period;
		Addr <=  "01000000011101";
		Trees_din <= x"02077504";
		wait for Clk_period;
		Addr <=  "01000000011110";
		Trees_din <= x"002140a9";
		wait for Clk_period;
		Addr <=  "01000000011111";
		Trees_din <= x"ffd540a9";
		wait for Clk_period;
		Addr <=  "01000000100000";
		Trees_din <= x"05f81704";
		wait for Clk_period;
		Addr <=  "01000000100001";
		Trees_din <= x"ffeb40a9";
		wait for Clk_period;
		Addr <=  "01000000100010";
		Trees_din <= x"006340a9";
		wait for Clk_period;
		Addr <=  "01000000100011";
		Trees_din <= x"0bf94704";
		wait for Clk_period;
		Addr <=  "01000000100100";
		Trees_din <= x"ffd640a9";
		wait for Clk_period;
		Addr <=  "01000000100101";
		Trees_din <= x"0b051f08";
		wait for Clk_period;
		Addr <=  "01000000100110";
		Trees_din <= x"0bfae404";
		wait for Clk_period;
		Addr <=  "01000000100111";
		Trees_din <= x"001840a9";
		wait for Clk_period;
		Addr <=  "01000000101000";
		Trees_din <= x"007e40a9";
		wait for Clk_period;
		Addr <=  "01000000101001";
		Trees_din <= x"fffa40a9";
		wait for Clk_period;
		Addr <=  "01000000101010";
		Trees_din <= x"000fd338";
		wait for Clk_period;
		Addr <=  "01000000101011";
		Trees_din <= x"03f63f0c";
		wait for Clk_period;
		Addr <=  "01000000101100";
		Trees_din <= x"11010d04";
		wait for Clk_period;
		Addr <=  "01000000101101";
		Trees_din <= x"001441c5";
		wait for Clk_period;
		Addr <=  "01000000101110";
		Trees_din <= x"04fa1604";
		wait for Clk_period;
		Addr <=  "01000000101111";
		Trees_din <= x"ff9341c5";
		wait for Clk_period;
		Addr <=  "01000000110000";
		Trees_din <= x"ffe541c5";
		wait for Clk_period;
		Addr <=  "01000000110001";
		Trees_din <= x"11fe7218";
		wait for Clk_period;
		Addr <=  "01000000110010";
		Trees_din <= x"0a030010";
		wait for Clk_period;
		Addr <=  "01000000110011";
		Trees_din <= x"09005408";
		wait for Clk_period;
		Addr <=  "01000000110100";
		Trees_din <= x"17000004";
		wait for Clk_period;
		Addr <=  "01000000110101";
		Trees_din <= x"005741c5";
		wait for Clk_period;
		Addr <=  "01000000110110";
		Trees_din <= x"001941c5";
		wait for Clk_period;
		Addr <=  "01000000110111";
		Trees_din <= x"09005a04";
		wait for Clk_period;
		Addr <=  "01000000111000";
		Trees_din <= x"ff9841c5";
		wait for Clk_period;
		Addr <=  "01000000111001";
		Trees_din <= x"003241c5";
		wait for Clk_period;
		Addr <=  "01000000111010";
		Trees_din <= x"10061504";
		wait for Clk_period;
		Addr <=  "01000000111011";
		Trees_din <= x"ff9441c5";
		wait for Clk_period;
		Addr <=  "01000000111100";
		Trees_din <= x"000e41c5";
		wait for Clk_period;
		Addr <=  "01000000111101";
		Trees_din <= x"0a044c0c";
		wait for Clk_period;
		Addr <=  "01000000111110";
		Trees_din <= x"0a03cc08";
		wait for Clk_period;
		Addr <=  "01000000111111";
		Trees_din <= x"09005d04";
		wait for Clk_period;
		Addr <=  "01000001000000";
		Trees_din <= x"fffd41c5";
		wait for Clk_period;
		Addr <=  "01000001000001";
		Trees_din <= x"004241c5";
		wait for Clk_period;
		Addr <=  "01000001000010";
		Trees_din <= x"ffb041c5";
		wait for Clk_period;
		Addr <=  "01000001000011";
		Trees_din <= x"13020c04";
		wait for Clk_period;
		Addr <=  "01000001000100";
		Trees_din <= x"006841c5";
		wait for Clk_period;
		Addr <=  "01000001000101";
		Trees_din <= x"000741c5";
		wait for Clk_period;
		Addr <=  "01000001000110";
		Trees_din <= x"17000424";
		wait for Clk_period;
		Addr <=  "01000001000111";
		Trees_din <= x"05f7e70c";
		wait for Clk_period;
		Addr <=  "01000001001000";
		Trees_din <= x"11027d08";
		wait for Clk_period;
		Addr <=  "01000001001001";
		Trees_din <= x"11016204";
		wait for Clk_period;
		Addr <=  "01000001001010";
		Trees_din <= x"002f41c5";
		wait for Clk_period;
		Addr <=  "01000001001011";
		Trees_din <= x"ffe841c5";
		wait for Clk_period;
		Addr <=  "01000001001100";
		Trees_din <= x"005c41c5";
		wait for Clk_period;
		Addr <=  "01000001001101";
		Trees_din <= x"09005108";
		wait for Clk_period;
		Addr <=  "01000001001110";
		Trees_din <= x"0b028804";
		wait for Clk_period;
		Addr <=  "01000001001111";
		Trees_din <= x"005a41c5";
		wait for Clk_period;
		Addr <=  "01000001010000";
		Trees_din <= x"ffea41c5";
		wait for Clk_period;
		Addr <=  "01000001010001";
		Trees_din <= x"07005808";
		wait for Clk_period;
		Addr <=  "01000001010010";
		Trees_din <= x"06f48004";
		wait for Clk_period;
		Addr <=  "01000001010011";
		Trees_din <= x"001a41c5";
		wait for Clk_period;
		Addr <=  "01000001010100";
		Trees_din <= x"ffad41c5";
		wait for Clk_period;
		Addr <=  "01000001010101";
		Trees_din <= x"0afc5304";
		wait for Clk_period;
		Addr <=  "01000001010110";
		Trees_din <= x"ffda41c5";
		wait for Clk_period;
		Addr <=  "01000001010111";
		Trees_din <= x"003f41c5";
		wait for Clk_period;
		Addr <=  "01000001011000";
		Trees_din <= x"0111441c";
		wait for Clk_period;
		Addr <=  "01000001011001";
		Trees_din <= x"1700690c";
		wait for Clk_period;
		Addr <=  "01000001011010";
		Trees_din <= x"07005b08";
		wait for Clk_period;
		Addr <=  "01000001011011";
		Trees_din <= x"10fa2804";
		wait for Clk_period;
		Addr <=  "01000001011100";
		Trees_din <= x"001c41c5";
		wait for Clk_period;
		Addr <=  "01000001011101";
		Trees_din <= x"008341c5";
		wait for Clk_period;
		Addr <=  "01000001011110";
		Trees_din <= x"ffee41c5";
		wait for Clk_period;
		Addr <=  "01000001011111";
		Trees_din <= x"1a00ce08";
		wait for Clk_period;
		Addr <=  "01000001100000";
		Trees_din <= x"08001e04";
		wait for Clk_period;
		Addr <=  "01000001100001";
		Trees_din <= x"004b41c5";
		wait for Clk_period;
		Addr <=  "01000001100010";
		Trees_din <= x"ffdb41c5";
		wait for Clk_period;
		Addr <=  "01000001100011";
		Trees_din <= x"1b003204";
		wait for Clk_period;
		Addr <=  "01000001100100";
		Trees_din <= x"ffec41c5";
		wait for Clk_period;
		Addr <=  "01000001100101";
		Trees_din <= x"007641c5";
		wait for Clk_period;
		Addr <=  "01000001100110";
		Trees_din <= x"0801b210";
		wait for Clk_period;
		Addr <=  "01000001100111";
		Trees_din <= x"00126b08";
		wait for Clk_period;
		Addr <=  "01000001101000";
		Trees_din <= x"05f92804";
		wait for Clk_period;
		Addr <=  "01000001101001";
		Trees_din <= x"ffa941c5";
		wait for Clk_period;
		Addr <=  "01000001101010";
		Trees_din <= x"001241c5";
		wait for Clk_period;
		Addr <=  "01000001101011";
		Trees_din <= x"11025d04";
		wait for Clk_period;
		Addr <=  "01000001101100";
		Trees_din <= x"001941c5";
		wait for Clk_period;
		Addr <=  "01000001101101";
		Trees_din <= x"005f41c5";
		wait for Clk_period;
		Addr <=  "01000001101110";
		Trees_din <= x"1101a204";
		wait for Clk_period;
		Addr <=  "01000001101111";
		Trees_din <= x"ffeb41c5";
		wait for Clk_period;
		Addr <=  "01000001110000";
		Trees_din <= x"ff9a41c5";
		wait for Clk_period;
		Addr <=  "01000001110001";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  2
        -----------
		Addr <=  "00000000000000";
		Trees_din <= x"03075d44";
		wait for Clk_period;
		Addr <=  "00000000000001";
		Trees_din <= x"03029118";
		wait for Clk_period;
		Addr <=  "00000000000010";
		Trees_din <= x"03004904";
		wait for Clk_period;
		Addr <=  "00000000000011";
		Trees_din <= x"ff4d0105";
		wait for Clk_period;
		Addr <=  "00000000000100";
		Trees_din <= x"07005e10";
		wait for Clk_period;
		Addr <=  "00000000000101";
		Trees_din <= x"0a034708";
		wait for Clk_period;
		Addr <=  "00000000000110";
		Trees_din <= x"0d03de04";
		wait for Clk_period;
		Addr <=  "00000000000111";
		Trees_din <= x"ff550105";
		wait for Clk_period;
		Addr <=  "00000000001000";
		Trees_din <= x"00270105";
		wait for Clk_period;
		Addr <=  "00000000001001";
		Trees_din <= x"0f003f04";
		wait for Clk_period;
		Addr <=  "00000000001010";
		Trees_din <= x"013c0105";
		wait for Clk_period;
		Addr <=  "00000000001011";
		Trees_din <= x"ff640105";
		wait for Clk_period;
		Addr <=  "00000000001100";
		Trees_din <= x"00590105";
		wait for Clk_period;
		Addr <=  "00000000001101";
		Trees_din <= x"06f54910";
		wait for Clk_period;
		Addr <=  "00000000001110";
		Trees_din <= x"1703a40c";
		wait for Clk_period;
		Addr <=  "00000000001111";
		Trees_din <= x"08000104";
		wait for Clk_period;
		Addr <=  "00000000010000";
		Trees_din <= x"00b20105";
		wait for Clk_period;
		Addr <=  "00000000010001";
		Trees_din <= x"01077d04";
		wait for Clk_period;
		Addr <=  "00000000010010";
		Trees_din <= x"ff530105";
		wait for Clk_period;
		Addr <=  "00000000010011";
		Trees_din <= x"00000105";
		wait for Clk_period;
		Addr <=  "00000000010100";
		Trees_din <= x"01290105";
		wait for Clk_period;
		Addr <=  "00000000010101";
		Trees_din <= x"04fc820c";
		wait for Clk_period;
		Addr <=  "00000000010110";
		Trees_din <= x"0104ee04";
		wait for Clk_period;
		Addr <=  "00000000010111";
		Trees_din <= x"ff590105";
		wait for Clk_period;
		Addr <=  "00000000011000";
		Trees_din <= x"0200f804";
		wait for Clk_period;
		Addr <=  "00000000011001";
		Trees_din <= x"ff9d0105";
		wait for Clk_period;
		Addr <=  "00000000011010";
		Trees_din <= x"010b0105";
		wait for Clk_period;
		Addr <=  "00000000011011";
		Trees_din <= x"00fba508";
		wait for Clk_period;
		Addr <=  "00000000011100";
		Trees_din <= x"01081404";
		wait for Clk_period;
		Addr <=  "00000000011101";
		Trees_din <= x"ff650105";
		wait for Clk_period;
		Addr <=  "00000000011110";
		Trees_din <= x"00270105";
		wait for Clk_period;
		Addr <=  "00000000011111";
		Trees_din <= x"07005a04";
		wait for Clk_period;
		Addr <=  "00000000100000";
		Trees_din <= x"007b0105";
		wait for Clk_period;
		Addr <=  "00000000100001";
		Trees_din <= x"02200105";
		wait for Clk_period;
		Addr <=  "00000000100010";
		Trees_din <= x"030a742c";
		wait for Clk_period;
		Addr <=  "00000000100011";
		Trees_din <= x"00fcaf18";
		wait for Clk_period;
		Addr <=  "00000000100100";
		Trees_din <= x"0c00e308";
		wait for Clk_period;
		Addr <=  "00000000100101";
		Trees_din <= x"01011d04";
		wait for Clk_period;
		Addr <=  "00000000100110";
		Trees_din <= x"ff7a0105";
		wait for Clk_period;
		Addr <=  "00000000100111";
		Trees_din <= x"00270105";
		wait for Clk_period;
		Addr <=  "00000000101000";
		Trees_din <= x"05fb7508";
		wait for Clk_period;
		Addr <=  "00000000101001";
		Trees_din <= x"0afc1404";
		wait for Clk_period;
		Addr <=  "00000000101010";
		Trees_din <= x"013c0105";
		wait for Clk_period;
		Addr <=  "00000000101011";
		Trees_din <= x"ffbb0105";
		wait for Clk_period;
		Addr <=  "00000000101100";
		Trees_din <= x"0100f904";
		wait for Clk_period;
		Addr <=  "00000000101101";
		Trees_din <= x"02a70105";
		wait for Clk_period;
		Addr <=  "00000000101110";
		Trees_din <= x"00b20105";
		wait for Clk_period;
		Addr <=  "00000000101111";
		Trees_din <= x"1202a108";
		wait for Clk_period;
		Addr <=  "00000000110000";
		Trees_din <= x"05fe5504";
		wait for Clk_period;
		Addr <=  "00000000110001";
		Trees_din <= x"035f0105";
		wait for Clk_period;
		Addr <=  "00000000110010";
		Trees_din <= x"01640105";
		wait for Clk_period;
		Addr <=  "00000000110011";
		Trees_din <= x"0f01f108";
		wait for Clk_period;
		Addr <=  "00000000110100";
		Trees_din <= x"06f52304";
		wait for Clk_period;
		Addr <=  "00000000110101";
		Trees_din <= x"00120105";
		wait for Clk_period;
		Addr <=  "00000000110110";
		Trees_din <= x"02030105";
		wait for Clk_period;
		Addr <=  "00000000110111";
		Trees_din <= x"ff9d0105";
		wait for Clk_period;
		Addr <=  "00000000111000";
		Trees_din <= x"0204ac10";
		wait for Clk_period;
		Addr <=  "00000000111001";
		Trees_din <= x"14001104";
		wait for Clk_period;
		Addr <=  "00000000111010";
		Trees_din <= x"00e20105";
		wait for Clk_period;
		Addr <=  "00000000111011";
		Trees_din <= x"05fec108";
		wait for Clk_period;
		Addr <=  "00000000111100";
		Trees_din <= x"06f3b404";
		wait for Clk_period;
		Addr <=  "00000000111101";
		Trees_din <= x"02720105";
		wait for Clk_period;
		Addr <=  "00000000111110";
		Trees_din <= x"03e30105";
		wait for Clk_period;
		Addr <=  "00000000111111";
		Trees_din <= x"013c0105";
		wait for Clk_period;
		Addr <=  "00000001000000";
		Trees_din <= x"00270105";
		wait for Clk_period;
		Addr <=  "00000001000001";
		Trees_din <= x"03063450";
		wait for Clk_period;
		Addr <=  "00000001000010";
		Trees_din <= x"03029118";
		wait for Clk_period;
		Addr <=  "00000001000011";
		Trees_din <= x"03004904";
		wait for Clk_period;
		Addr <=  "00000001000100";
		Trees_din <= x"ff540211";
		wait for Clk_period;
		Addr <=  "00000001000101";
		Trees_din <= x"07005e10";
		wait for Clk_period;
		Addr <=  "00000001000110";
		Trees_din <= x"1005e408";
		wait for Clk_period;
		Addr <=  "00000001000111";
		Trees_din <= x"05015d04";
		wait for Clk_period;
		Addr <=  "00000001001000";
		Trees_din <= x"ff600211";
		wait for Clk_period;
		Addr <=  "00000001001001";
		Trees_din <= x"00280211";
		wait for Clk_period;
		Addr <=  "00000001001010";
		Trees_din <= x"14016904";
		wait for Clk_period;
		Addr <=  "00000001001011";
		Trees_din <= x"00d10211";
		wait for Clk_period;
		Addr <=  "00000001001100";
		Trees_din <= x"ff840211";
		wait for Clk_period;
		Addr <=  "00000001001101";
		Trees_din <= x"00580211";
		wait for Clk_period;
		Addr <=  "00000001001110";
		Trees_din <= x"0c016e1c";
		wait for Clk_period;
		Addr <=  "00000001001111";
		Trees_din <= x"1900a810";
		wait for Clk_period;
		Addr <=  "00000001010000";
		Trees_din <= x"1b004808";
		wait for Clk_period;
		Addr <=  "00000001010001";
		Trees_din <= x"0c00e904";
		wait for Clk_period;
		Addr <=  "00000001010010";
		Trees_din <= x"ff760211";
		wait for Clk_period;
		Addr <=  "00000001010011";
		Trees_din <= x"00400211";
		wait for Clk_period;
		Addr <=  "00000001010100";
		Trees_din <= x"0101ee04";
		wait for Clk_period;
		Addr <=  "00000001010101";
		Trees_din <= x"ffc40211";
		wait for Clk_period;
		Addr <=  "00000001010110";
		Trees_din <= x"01ce0211";
		wait for Clk_period;
		Addr <=  "00000001010111";
		Trees_din <= x"1b002e08";
		wait for Clk_period;
		Addr <=  "00000001011000";
		Trees_din <= x"1500a704";
		wait for Clk_period;
		Addr <=  "00000001011001";
		Trees_din <= x"ff9d0211";
		wait for Clk_period;
		Addr <=  "00000001011010";
		Trees_din <= x"00cd0211";
		wait for Clk_period;
		Addr <=  "00000001011011";
		Trees_din <= x"01e40211";
		wait for Clk_period;
		Addr <=  "00000001011100";
		Trees_din <= x"2004000c";
		wait for Clk_period;
		Addr <=  "00000001011101";
		Trees_din <= x"13fec408";
		wait for Clk_period;
		Addr <=  "00000001011110";
		Trees_din <= x"04016e04";
		wait for Clk_period;
		Addr <=  "00000001011111";
		Trees_din <= x"00050211";
		wait for Clk_period;
		Addr <=  "00000001100000";
		Trees_din <= x"01b80211";
		wait for Clk_period;
		Addr <=  "00000001100001";
		Trees_din <= x"ff820211";
		wait for Clk_period;
		Addr <=  "00000001100010";
		Trees_din <= x"0305c708";
		wait for Clk_period;
		Addr <=  "00000001100011";
		Trees_din <= x"12040104";
		wait for Clk_period;
		Addr <=  "00000001100100";
		Trees_din <= x"ff6d0211";
		wait for Clk_period;
		Addr <=  "00000001100101";
		Trees_din <= x"00370211";
		wait for Clk_period;
		Addr <=  "00000001100110";
		Trees_din <= x"10045104";
		wait for Clk_period;
		Addr <=  "00000001100111";
		Trees_din <= x"ff800211";
		wait for Clk_period;
		Addr <=  "00000001101000";
		Trees_din <= x"01320211";
		wait for Clk_period;
		Addr <=  "00000001101001";
		Trees_din <= x"0307f520";
		wait for Clk_period;
		Addr <=  "00000001101010";
		Trees_din <= x"05f92808";
		wait for Clk_period;
		Addr <=  "00000001101011";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00000001101100";
		Trees_din <= x"003b0211";
		wait for Clk_period;
		Addr <=  "00000001101101";
		Trees_din <= x"ff700211";
		wait for Clk_period;
		Addr <=  "00000001101110";
		Trees_din <= x"17000b0c";
		wait for Clk_period;
		Addr <=  "00000001101111";
		Trees_din <= x"0c01c808";
		wait for Clk_period;
		Addr <=  "00000001110000";
		Trees_din <= x"0400ad04";
		wait for Clk_period;
		Addr <=  "00000001110001";
		Trees_din <= x"013d0211";
		wait for Clk_period;
		Addr <=  "00000001110010";
		Trees_din <= x"fff70211";
		wait for Clk_period;
		Addr <=  "00000001110011";
		Trees_din <= x"ff780211";
		wait for Clk_period;
		Addr <=  "00000001110100";
		Trees_din <= x"18003304";
		wait for Clk_period;
		Addr <=  "00000001110101";
		Trees_din <= x"ff8c0211";
		wait for Clk_period;
		Addr <=  "00000001110110";
		Trees_din <= x"0202c504";
		wait for Clk_period;
		Addr <=  "00000001110111";
		Trees_din <= x"01900211";
		wait for Clk_period;
		Addr <=  "00000001111000";
		Trees_din <= x"00060211";
		wait for Clk_period;
		Addr <=  "00000001111001";
		Trees_din <= x"0204ac10";
		wait for Clk_period;
		Addr <=  "00000001111010";
		Trees_din <= x"0803ed0c";
		wait for Clk_period;
		Addr <=  "00000001111011";
		Trees_din <= x"00050808";
		wait for Clk_period;
		Addr <=  "00000001111100";
		Trees_din <= x"1a00a104";
		wait for Clk_period;
		Addr <=  "00000001111101";
		Trees_din <= x"011c0211";
		wait for Clk_period;
		Addr <=  "00000001111110";
		Trees_din <= x"019e0211";
		wait for Clk_period;
		Addr <=  "00000001111111";
		Trees_din <= x"006a0211";
		wait for Clk_period;
		Addr <=  "00000010000000";
		Trees_din <= x"00260211";
		wait for Clk_period;
		Addr <=  "00000010000001";
		Trees_din <= x"0effa704";
		wait for Clk_period;
		Addr <=  "00000010000010";
		Trees_din <= x"00bb0211";
		wait for Clk_period;
		Addr <=  "00000010000011";
		Trees_din <= x"ff8b0211";
		wait for Clk_period;
		Addr <=  "00000010000100";
		Trees_din <= x"03063448";
		wait for Clk_period;
		Addr <=  "00000010000101";
		Trees_din <= x"0302911c";
		wait for Clk_period;
		Addr <=  "00000010000110";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00000010000111";
		Trees_din <= x"ff580325";
		wait for Clk_period;
		Addr <=  "00000010001000";
		Trees_din <= x"07005e10";
		wait for Clk_period;
		Addr <=  "00000010001001";
		Trees_din <= x"08000908";
		wait for Clk_period;
		Addr <=  "00000010001010";
		Trees_din <= x"0000af04";
		wait for Clk_period;
		Addr <=  "00000010001011";
		Trees_din <= x"00640325";
		wait for Clk_period;
		Addr <=  "00000010001100";
		Trees_din <= x"ff770325";
		wait for Clk_period;
		Addr <=  "00000010001101";
		Trees_din <= x"1005e404";
		wait for Clk_period;
		Addr <=  "00000010001110";
		Trees_din <= x"ff5f0325";
		wait for Clk_period;
		Addr <=  "00000010001111";
		Trees_din <= x"ffc40325";
		wait for Clk_period;
		Addr <=  "00000010010000";
		Trees_din <= x"0efebe04";
		wait for Clk_period;
		Addr <=  "00000010010001";
		Trees_din <= x"01030325";
		wait for Clk_period;
		Addr <=  "00000010010010";
		Trees_din <= x"ff820325";
		wait for Clk_period;
		Addr <=  "00000010010011";
		Trees_din <= x"0c016e14";
		wait for Clk_period;
		Addr <=  "00000010010100";
		Trees_din <= x"00fae404";
		wait for Clk_period;
		Addr <=  "00000010010101";
		Trees_din <= x"ff6f0325";
		wait for Clk_period;
		Addr <=  "00000010010110";
		Trees_din <= x"0101d108";
		wait for Clk_period;
		Addr <=  "00000010010111";
		Trees_din <= x"1c002e04";
		wait for Clk_period;
		Addr <=  "00000010011000";
		Trees_din <= x"01150325";
		wait for Clk_period;
		Addr <=  "00000010011001";
		Trees_din <= x"ff960325";
		wait for Clk_period;
		Addr <=  "00000010011010";
		Trees_din <= x"1b002e04";
		wait for Clk_period;
		Addr <=  "00000010011011";
		Trees_din <= x"ff980325";
		wait for Clk_period;
		Addr <=  "00000010011100";
		Trees_din <= x"01270325";
		wait for Clk_period;
		Addr <=  "00000010011101";
		Trees_din <= x"2004000c";
		wait for Clk_period;
		Addr <=  "00000010011110";
		Trees_din <= x"13fec408";
		wait for Clk_period;
		Addr <=  "00000010011111";
		Trees_din <= x"0f017804";
		wait for Clk_period;
		Addr <=  "00000010100000";
		Trees_din <= x"01490325";
		wait for Clk_period;
		Addr <=  "00000010100001";
		Trees_din <= x"fff40325";
		wait for Clk_period;
		Addr <=  "00000010100010";
		Trees_din <= x"ff890325";
		wait for Clk_period;
		Addr <=  "00000010100011";
		Trees_din <= x"0a015608";
		wait for Clk_period;
		Addr <=  "00000010100100";
		Trees_din <= x"13fd5204";
		wait for Clk_period;
		Addr <=  "00000010100101";
		Trees_din <= x"009d0325";
		wait for Clk_period;
		Addr <=  "00000010100110";
		Trees_din <= x"ffb00325";
		wait for Clk_period;
		Addr <=  "00000010100111";
		Trees_din <= x"ff5b0325";
		wait for Clk_period;
		Addr <=  "00000010101000";
		Trees_din <= x"0308a924";
		wait for Clk_period;
		Addr <=  "00000010101001";
		Trees_din <= x"05f86604";
		wait for Clk_period;
		Addr <=  "00000010101010";
		Trees_din <= x"ff7c0325";
		wait for Clk_period;
		Addr <=  "00000010101011";
		Trees_din <= x"07005910";
		wait for Clk_period;
		Addr <=  "00000010101100";
		Trees_din <= x"0bfacb08";
		wait for Clk_period;
		Addr <=  "00000010101101";
		Trees_din <= x"0306c204";
		wait for Clk_period;
		Addr <=  "00000010101110";
		Trees_din <= x"009a0325";
		wait for Clk_period;
		Addr <=  "00000010101111";
		Trees_din <= x"ff640325";
		wait for Clk_period;
		Addr <=  "00000010110000";
		Trees_din <= x"1d003d04";
		wait for Clk_period;
		Addr <=  "00000010110001";
		Trees_din <= x"01280325";
		wait for Clk_period;
		Addr <=  "00000010110010";
		Trees_din <= x"00200325";
		wait for Clk_period;
		Addr <=  "00000010110011";
		Trees_din <= x"02016008";
		wait for Clk_period;
		Addr <=  "00000010110100";
		Trees_din <= x"01fcbe04";
		wait for Clk_period;
		Addr <=  "00000010110101";
		Trees_din <= x"001b0325";
		wait for Clk_period;
		Addr <=  "00000010110110";
		Trees_din <= x"01790325";
		wait for Clk_period;
		Addr <=  "00000010110111";
		Trees_din <= x"12013204";
		wait for Clk_period;
		Addr <=  "00000010111000";
		Trees_din <= x"00bd0325";
		wait for Clk_period;
		Addr <=  "00000010111001";
		Trees_din <= x"ff900325";
		wait for Clk_period;
		Addr <=  "00000010111010";
		Trees_din <= x"0204ac18";
		wait for Clk_period;
		Addr <=  "00000010111011";
		Trees_din <= x"0c00290c";
		wait for Clk_period;
		Addr <=  "00000010111100";
		Trees_din <= x"030bbf04";
		wait for Clk_period;
		Addr <=  "00000010111101";
		Trees_din <= x"ff790325";
		wait for Clk_period;
		Addr <=  "00000010111110";
		Trees_din <= x"05fa0504";
		wait for Clk_period;
		Addr <=  "00000010111111";
		Trees_din <= x"00420325";
		wait for Clk_period;
		Addr <=  "00000011000000";
		Trees_din <= x"01240325";
		wait for Clk_period;
		Addr <=  "00000011000001";
		Trees_din <= x"1f003208";
		wait for Clk_period;
		Addr <=  "00000011000010";
		Trees_din <= x"10f72e04";
		wait for Clk_period;
		Addr <=  "00000011000011";
		Trees_din <= x"00910325";
		wait for Clk_period;
		Addr <=  "00000011000100";
		Trees_din <= x"01280325";
		wait for Clk_period;
		Addr <=  "00000011000101";
		Trees_din <= x"003b0325";
		wait for Clk_period;
		Addr <=  "00000011000110";
		Trees_din <= x"11ff9e04";
		wait for Clk_period;
		Addr <=  "00000011000111";
		Trees_din <= x"00c80325";
		wait for Clk_period;
		Addr <=  "00000011001000";
		Trees_din <= x"ff8a0325";
		wait for Clk_period;
		Addr <=  "00000011001001";
		Trees_din <= x"0304d348";
		wait for Clk_period;
		Addr <=  "00000011001010";
		Trees_din <= x"0301f918";
		wait for Clk_period;
		Addr <=  "00000011001011";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00000011001100";
		Trees_din <= x"ff5c0459";
		wait for Clk_period;
		Addr <=  "00000011001101";
		Trees_din <= x"1f001410";
		wait for Clk_period;
		Addr <=  "00000011001110";
		Trees_din <= x"07005e08";
		wait for Clk_period;
		Addr <=  "00000011001111";
		Trees_din <= x"11048e04";
		wait for Clk_period;
		Addr <=  "00000011010000";
		Trees_din <= x"ff640459";
		wait for Clk_period;
		Addr <=  "00000011010001";
		Trees_din <= x"fff80459";
		wait for Clk_period;
		Addr <=  "00000011010010";
		Trees_din <= x"0efe7004";
		wait for Clk_period;
		Addr <=  "00000011010011";
		Trees_din <= x"00c20459";
		wait for Clk_period;
		Addr <=  "00000011010100";
		Trees_din <= x"ff960459";
		wait for Clk_period;
		Addr <=  "00000011010101";
		Trees_din <= x"00730459";
		wait for Clk_period;
		Addr <=  "00000011010110";
		Trees_din <= x"0e001a1c";
		wait for Clk_period;
		Addr <=  "00000011010111";
		Trees_din <= x"0f008c10";
		wait for Clk_period;
		Addr <=  "00000011011000";
		Trees_din <= x"0303cb08";
		wait for Clk_period;
		Addr <=  "00000011011001";
		Trees_din <= x"0204e504";
		wait for Clk_period;
		Addr <=  "00000011011010";
		Trees_din <= x"01490459";
		wait for Clk_period;
		Addr <=  "00000011011011";
		Trees_din <= x"ffa70459";
		wait for Clk_period;
		Addr <=  "00000011011100";
		Trees_din <= x"01ffc504";
		wait for Clk_period;
		Addr <=  "00000011011101";
		Trees_din <= x"00300459";
		wait for Clk_period;
		Addr <=  "00000011011110";
		Trees_din <= x"ff8e0459";
		wait for Clk_period;
		Addr <=  "00000011011111";
		Trees_din <= x"07005004";
		wait for Clk_period;
		Addr <=  "00000011100000";
		Trees_din <= x"011e0459";
		wait for Clk_period;
		Addr <=  "00000011100001";
		Trees_din <= x"10028004";
		wait for Clk_period;
		Addr <=  "00000011100010";
		Trees_din <= x"00030459";
		wait for Clk_period;
		Addr <=  "00000011100011";
		Trees_din <= x"ff640459";
		wait for Clk_period;
		Addr <=  "00000011100100";
		Trees_din <= x"08000308";
		wait for Clk_period;
		Addr <=  "00000011100101";
		Trees_din <= x"01042f04";
		wait for Clk_period;
		Addr <=  "00000011100110";
		Trees_din <= x"ffa20459";
		wait for Clk_period;
		Addr <=  "00000011100111";
		Trees_din <= x"00f60459";
		wait for Clk_period;
		Addr <=  "00000011101000";
		Trees_din <= x"07004804";
		wait for Clk_period;
		Addr <=  "00000011101001";
		Trees_din <= x"00880459";
		wait for Clk_period;
		Addr <=  "00000011101010";
		Trees_din <= x"05ff6b04";
		wait for Clk_period;
		Addr <=  "00000011101011";
		Trees_din <= x"ff640459";
		wait for Clk_period;
		Addr <=  "00000011101100";
		Trees_din <= x"00430459";
		wait for Clk_period;
		Addr <=  "00000011101101";
		Trees_din <= x"0307f534";
		wait for Clk_period;
		Addr <=  "00000011101110";
		Trees_din <= x"0800f020";
		wait for Clk_period;
		Addr <=  "00000011101111";
		Trees_din <= x"08007b10";
		wait for Clk_period;
		Addr <=  "00000011110000";
		Trees_din <= x"06f5d008";
		wait for Clk_period;
		Addr <=  "00000011110001";
		Trees_din <= x"0b04f204";
		wait for Clk_period;
		Addr <=  "00000011110010";
		Trees_din <= x"ff6e0459";
		wait for Clk_period;
		Addr <=  "00000011110011";
		Trees_din <= x"00150459";
		wait for Clk_period;
		Addr <=  "00000011110100";
		Trees_din <= x"14007a04";
		wait for Clk_period;
		Addr <=  "00000011110101";
		Trees_din <= x"ffc60459";
		wait for Clk_period;
		Addr <=  "00000011110110";
		Trees_din <= x"00bf0459";
		wait for Clk_period;
		Addr <=  "00000011110111";
		Trees_din <= x"0f017808";
		wait for Clk_period;
		Addr <=  "00000011111000";
		Trees_din <= x"05f9e904";
		wait for Clk_period;
		Addr <=  "00000011111001";
		Trees_din <= x"00670459";
		wait for Clk_period;
		Addr <=  "00000011111010";
		Trees_din <= x"01a10459";
		wait for Clk_period;
		Addr <=  "00000011111011";
		Trees_din <= x"11006c04";
		wait for Clk_period;
		Addr <=  "00000011111100";
		Trees_din <= x"00d30459";
		wait for Clk_period;
		Addr <=  "00000011111101";
		Trees_din <= x"ff8d0459";
		wait for Clk_period;
		Addr <=  "00000011111110";
		Trees_din <= x"08020104";
		wait for Clk_period;
		Addr <=  "00000011111111";
		Trees_din <= x"ff5c0459";
		wait for Clk_period;
		Addr <=  "00000100000000";
		Trees_din <= x"16035e08";
		wait for Clk_period;
		Addr <=  "00000100000001";
		Trees_din <= x"10059d04";
		wait for Clk_period;
		Addr <=  "00000100000010";
		Trees_din <= x"ff7d0459";
		wait for Clk_period;
		Addr <=  "00000100000011";
		Trees_din <= x"00f90459";
		wait for Clk_period;
		Addr <=  "00000100000100";
		Trees_din <= x"0afc3704";
		wait for Clk_period;
		Addr <=  "00000100000101";
		Trees_din <= x"fffd0459";
		wait for Clk_period;
		Addr <=  "00000100000110";
		Trees_din <= x"00f40459";
		wait for Clk_period;
		Addr <=  "00000100000111";
		Trees_din <= x"0410f71c";
		wait for Clk_period;
		Addr <=  "00000100001000";
		Trees_din <= x"030da80c";
		wait for Clk_period;
		Addr <=  "00000100001001";
		Trees_din <= x"18005508";
		wait for Clk_period;
		Addr <=  "00000100001010";
		Trees_din <= x"1500b104";
		wait for Clk_period;
		Addr <=  "00000100001011";
		Trees_din <= x"00c60459";
		wait for Clk_period;
		Addr <=  "00000100001100";
		Trees_din <= x"ffb90459";
		wait for Clk_period;
		Addr <=  "00000100001101";
		Trees_din <= x"ff790459";
		wait for Clk_period;
		Addr <=  "00000100001110";
		Trees_din <= x"1104d508";
		wait for Clk_period;
		Addr <=  "00000100001111";
		Trees_din <= x"05f54504";
		wait for Clk_period;
		Addr <=  "00000100010000";
		Trees_din <= x"00480459";
		wait for Clk_period;
		Addr <=  "00000100010001";
		Trees_din <= x"01050459";
		wait for Clk_period;
		Addr <=  "00000100010010";
		Trees_din <= x"07005604";
		wait for Clk_period;
		Addr <=  "00000100010011";
		Trees_din <= x"00a90459";
		wait for Clk_period;
		Addr <=  "00000100010100";
		Trees_din <= x"ffbd0459";
		wait for Clk_period;
		Addr <=  "00000100010101";
		Trees_din <= x"ff8f0459";
		wait for Clk_period;
		Addr <=  "00000100010110";
		Trees_din <= x"0304d348";
		wait for Clk_period;
		Addr <=  "00000100010111";
		Trees_din <= x"0301f91c";
		wait for Clk_period;
		Addr <=  "00000100011000";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00000100011001";
		Trees_din <= x"ff5e0585";
		wait for Clk_period;
		Addr <=  "00000100011010";
		Trees_din <= x"07005e10";
		wait for Clk_period;
		Addr <=  "00000100011011";
		Trees_din <= x"08000908";
		wait for Clk_period;
		Addr <=  "00000100011100";
		Trees_din <= x"0bfad604";
		wait for Clk_period;
		Addr <=  "00000100011101";
		Trees_din <= x"00a40585";
		wait for Clk_period;
		Addr <=  "00000100011110";
		Trees_din <= x"ff850585";
		wait for Clk_period;
		Addr <=  "00000100011111";
		Trees_din <= x"1b002d04";
		wait for Clk_period;
		Addr <=  "00000100100000";
		Trees_din <= x"ffb70585";
		wait for Clk_period;
		Addr <=  "00000100100001";
		Trees_din <= x"ff5f0585";
		wait for Clk_period;
		Addr <=  "00000100100010";
		Trees_din <= x"0202b804";
		wait for Clk_period;
		Addr <=  "00000100100011";
		Trees_din <= x"ff8f0585";
		wait for Clk_period;
		Addr <=  "00000100100100";
		Trees_din <= x"00da0585";
		wait for Clk_period;
		Addr <=  "00000100100101";
		Trees_din <= x"0efe9614";
		wait for Clk_period;
		Addr <=  "00000100100110";
		Trees_din <= x"06f40d04";
		wait for Clk_period;
		Addr <=  "00000100100111";
		Trees_din <= x"ff7f0585";
		wait for Clk_period;
		Addr <=  "00000100101000";
		Trees_din <= x"09005508";
		wait for Clk_period;
		Addr <=  "00000100101001";
		Trees_din <= x"1500a504";
		wait for Clk_period;
		Addr <=  "00000100101010";
		Trees_din <= x"01180585";
		wait for Clk_period;
		Addr <=  "00000100101011";
		Trees_din <= x"00060585";
		wait for Clk_period;
		Addr <=  "00000100101100";
		Trees_din <= x"0c032604";
		wait for Clk_period;
		Addr <=  "00000100101101";
		Trees_din <= x"ff7d0585";
		wait for Clk_period;
		Addr <=  "00000100101110";
		Trees_din <= x"00790585";
		wait for Clk_period;
		Addr <=  "00000100101111";
		Trees_din <= x"08000308";
		wait for Clk_period;
		Addr <=  "00000100110000";
		Trees_din <= x"01042f04";
		wait for Clk_period;
		Addr <=  "00000100110001";
		Trees_din <= x"ffa70585";
		wait for Clk_period;
		Addr <=  "00000100110010";
		Trees_din <= x"00e50585";
		wait for Clk_period;
		Addr <=  "00000100110011";
		Trees_din <= x"08026908";
		wait for Clk_period;
		Addr <=  "00000100110100";
		Trees_din <= x"1703e904";
		wait for Clk_period;
		Addr <=  "00000100110101";
		Trees_din <= x"ff660585";
		wait for Clk_period;
		Addr <=  "00000100110110";
		Trees_din <= x"00530585";
		wait for Clk_period;
		Addr <=  "00000100110111";
		Trees_din <= x"18004004";
		wait for Clk_period;
		Addr <=  "00000100111000";
		Trees_din <= x"ffad0585";
		wait for Clk_period;
		Addr <=  "00000100111001";
		Trees_din <= x"012d0585";
		wait for Clk_period;
		Addr <=  "00000100111010";
		Trees_din <= x"0308a930";
		wait for Clk_period;
		Addr <=  "00000100111011";
		Trees_din <= x"0800f01c";
		wait for Clk_period;
		Addr <=  "00000100111100";
		Trees_din <= x"08007b10";
		wait for Clk_period;
		Addr <=  "00000100111101";
		Trees_din <= x"09005708";
		wait for Clk_period;
		Addr <=  "00000100111110";
		Trees_din <= x"0c028204";
		wait for Clk_period;
		Addr <=  "00000100111111";
		Trees_din <= x"ffb60585";
		wait for Clk_period;
		Addr <=  "00000101000000";
		Trees_din <= x"00940585";
		wait for Clk_period;
		Addr <=  "00000101000001";
		Trees_din <= x"0f000704";
		wait for Clk_period;
		Addr <=  "00000101000010";
		Trees_din <= x"ffa40585";
		wait for Clk_period;
		Addr <=  "00000101000011";
		Trees_din <= x"00b40585";
		wait for Clk_period;
		Addr <=  "00000101000100";
		Trees_din <= x"05f86604";
		wait for Clk_period;
		Addr <=  "00000101000101";
		Trees_din <= x"ff9e0585";
		wait for Clk_period;
		Addr <=  "00000101000110";
		Trees_din <= x"16005604";
		wait for Clk_period;
		Addr <=  "00000101000111";
		Trees_din <= x"003b0585";
		wait for Clk_period;
		Addr <=  "00000101001000";
		Trees_din <= x"01330585";
		wait for Clk_period;
		Addr <=  "00000101001001";
		Trees_din <= x"0305c704";
		wait for Clk_period;
		Addr <=  "00000101001010";
		Trees_din <= x"ff6f0585";
		wait for Clk_period;
		Addr <=  "00000101001011";
		Trees_din <= x"00fe7b08";
		wait for Clk_period;
		Addr <=  "00000101001100";
		Trees_din <= x"1900aa04";
		wait for Clk_period;
		Addr <=  "00000101001101";
		Trees_din <= x"ff9e0585";
		wait for Clk_period;
		Addr <=  "00000101001110";
		Trees_din <= x"00710585";
		wait for Clk_period;
		Addr <=  "00000101001111";
		Trees_din <= x"1c003604";
		wait for Clk_period;
		Addr <=  "00000101010000";
		Trees_din <= x"00920585";
		wait for Clk_period;
		Addr <=  "00000101010001";
		Trees_din <= x"ff840585";
		wait for Clk_period;
		Addr <=  "00000101010010";
		Trees_din <= x"0204ac18";
		wait for Clk_period;
		Addr <=  "00000101010011";
		Trees_din <= x"06f0dc08";
		wait for Clk_period;
		Addr <=  "00000101010100";
		Trees_din <= x"02014b04";
		wait for Clk_period;
		Addr <=  "00000101010101";
		Trees_din <= x"ff7d0585";
		wait for Clk_period;
		Addr <=  "00000101010110";
		Trees_din <= x"006f0585";
		wait for Clk_period;
		Addr <=  "00000101010111";
		Trees_din <= x"030da808";
		wait for Clk_period;
		Addr <=  "00000101011000";
		Trees_din <= x"14001104";
		wait for Clk_period;
		Addr <=  "00000101011001";
		Trees_din <= x"ff970585";
		wait for Clk_period;
		Addr <=  "00000101011010";
		Trees_din <= x"00a80585";
		wait for Clk_period;
		Addr <=  "00000101011011";
		Trees_din <= x"0c03e204";
		wait for Clk_period;
		Addr <=  "00000101011100";
		Trees_din <= x"00db0585";
		wait for Clk_period;
		Addr <=  "00000101011101";
		Trees_din <= x"00320585";
		wait for Clk_period;
		Addr <=  "00000101011110";
		Trees_din <= x"11ff9e04";
		wait for Clk_period;
		Addr <=  "00000101011111";
		Trees_din <= x"00920585";
		wait for Clk_period;
		Addr <=  "00000101100000";
		Trees_din <= x"ff890585";
		wait for Clk_period;
		Addr <=  "00000101100001";
		Trees_din <= x"0304d344";
		wait for Clk_period;
		Addr <=  "00000101100010";
		Trees_din <= x"0301f918";
		wait for Clk_period;
		Addr <=  "00000101100011";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00000101100100";
		Trees_din <= x"ff600689";
		wait for Clk_period;
		Addr <=  "00000101100101";
		Trees_din <= x"1f001410";
		wait for Clk_period;
		Addr <=  "00000101100110";
		Trees_din <= x"07005e08";
		wait for Clk_period;
		Addr <=  "00000101100111";
		Trees_din <= x"11048e04";
		wait for Clk_period;
		Addr <=  "00000101101000";
		Trees_din <= x"ff6d0689";
		wait for Clk_period;
		Addr <=  "00000101101001";
		Trees_din <= x"00100689";
		wait for Clk_period;
		Addr <=  "00000101101010";
		Trees_din <= x"0efe7004";
		wait for Clk_period;
		Addr <=  "00000101101011";
		Trees_din <= x"00ac0689";
		wait for Clk_period;
		Addr <=  "00000101101100";
		Trees_din <= x"ff9a0689";
		wait for Clk_period;
		Addr <=  "00000101101101";
		Trees_din <= x"00780689";
		wait for Clk_period;
		Addr <=  "00000101101110";
		Trees_din <= x"12fe8d10";
		wait for Clk_period;
		Addr <=  "00000101101111";
		Trees_din <= x"12fe440c";
		wait for Clk_period;
		Addr <=  "00000101110000";
		Trees_din <= x"0a036d04";
		wait for Clk_period;
		Addr <=  "00000101110001";
		Trees_din <= x"ff770689";
		wait for Clk_period;
		Addr <=  "00000101110010";
		Trees_din <= x"0a046704";
		wait for Clk_period;
		Addr <=  "00000101110011";
		Trees_din <= x"00c30689";
		wait for Clk_period;
		Addr <=  "00000101110100";
		Trees_din <= x"ff9b0689";
		wait for Clk_period;
		Addr <=  "00000101110101";
		Trees_din <= x"012a0689";
		wait for Clk_period;
		Addr <=  "00000101110110";
		Trees_din <= x"05ff6b10";
		wait for Clk_period;
		Addr <=  "00000101110111";
		Trees_din <= x"1f000008";
		wait for Clk_period;
		Addr <=  "00000101111000";
		Trees_din <= x"08000304";
		wait for Clk_period;
		Addr <=  "00000101111001";
		Trees_din <= x"003c0689";
		wait for Clk_period;
		Addr <=  "00000101111010";
		Trees_din <= x"ff7d0689";
		wait for Clk_period;
		Addr <=  "00000101111011";
		Trees_din <= x"0d003904";
		wait for Clk_period;
		Addr <=  "00000101111100";
		Trees_din <= x"00b70689";
		wait for Clk_period;
		Addr <=  "00000101111101";
		Trees_din <= x"ffc50689";
		wait for Clk_period;
		Addr <=  "00000101111110";
		Trees_din <= x"05ffbc04";
		wait for Clk_period;
		Addr <=  "00000101111111";
		Trees_din <= x"01170689";
		wait for Clk_period;
		Addr <=  "00000110000000";
		Trees_din <= x"0f012e04";
		wait for Clk_period;
		Addr <=  "00000110000001";
		Trees_din <= x"ff9d0689";
		wait for Clk_period;
		Addr <=  "00000110000010";
		Trees_din <= x"00240689";
		wait for Clk_period;
		Addr <=  "00000110000011";
		Trees_din <= x"030bbf1c";
		wait for Clk_period;
		Addr <=  "00000110000100";
		Trees_din <= x"02053814";
		wait for Clk_period;
		Addr <=  "00000110000101";
		Trees_din <= x"0c002904";
		wait for Clk_period;
		Addr <=  "00000110000110";
		Trees_din <= x"ff670689";
		wait for Clk_period;
		Addr <=  "00000110000111";
		Trees_din <= x"07005908";
		wait for Clk_period;
		Addr <=  "00000110001000";
		Trees_din <= x"1e006b04";
		wait for Clk_period;
		Addr <=  "00000110001001";
		Trees_din <= x"006a0689";
		wait for Clk_period;
		Addr <=  "00000110001010";
		Trees_din <= x"fff70689";
		wait for Clk_period;
		Addr <=  "00000110001011";
		Trees_din <= x"00fa2404";
		wait for Clk_period;
		Addr <=  "00000110001100";
		Trees_din <= x"ffe40689";
		wait for Clk_period;
		Addr <=  "00000110001101";
		Trees_din <= x"00b50689";
		wait for Clk_period;
		Addr <=  "00000110001110";
		Trees_din <= x"09005904";
		wait for Clk_period;
		Addr <=  "00000110001111";
		Trees_din <= x"ff6e0689";
		wait for Clk_period;
		Addr <=  "00000110010000";
		Trees_din <= x"00040689";
		wait for Clk_period;
		Addr <=  "00000110010001";
		Trees_din <= x"040a4a14";
		wait for Clk_period;
		Addr <=  "00000110010010";
		Trees_din <= x"05fec110";
		wait for Clk_period;
		Addr <=  "00000110010011";
		Trees_din <= x"05f54508";
		wait for Clk_period;
		Addr <=  "00000110010100";
		Trees_din <= x"0b028704";
		wait for Clk_period;
		Addr <=  "00000110010101";
		Trees_din <= x"00890689";
		wait for Clk_period;
		Addr <=  "00000110010110";
		Trees_din <= x"ff880689";
		wait for Clk_period;
		Addr <=  "00000110010111";
		Trees_din <= x"1104d504";
		wait for Clk_period;
		Addr <=  "00000110011000";
		Trees_din <= x"00c70689";
		wait for Clk_period;
		Addr <=  "00000110011001";
		Trees_din <= x"003a0689";
		wait for Clk_period;
		Addr <=  "00000110011010";
		Trees_din <= x"fff90689";
		wait for Clk_period;
		Addr <=  "00000110011011";
		Trees_din <= x"0f012b0c";
		wait for Clk_period;
		Addr <=  "00000110011100";
		Trees_din <= x"15009b08";
		wait for Clk_period;
		Addr <=  "00000110011101";
		Trees_din <= x"19009704";
		wait for Clk_period;
		Addr <=  "00000110011110";
		Trees_din <= x"fffb0689";
		wait for Clk_period;
		Addr <=  "00000110011111";
		Trees_din <= x"ff3d0689";
		wait for Clk_period;
		Addr <=  "00000110100000";
		Trees_din <= x"00890689";
		wait for Clk_period;
		Addr <=  "00000110100001";
		Trees_din <= x"00be0689";
		wait for Clk_period;
		Addr <=  "00000110100010";
		Trees_din <= x"03029128";
		wait for Clk_period;
		Addr <=  "00000110100011";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00000110100100";
		Trees_din <= x"ff620765";
		wait for Clk_period;
		Addr <=  "00000110100101";
		Trees_din <= x"07005e1c";
		wait for Clk_period;
		Addr <=  "00000110100110";
		Trees_din <= x"0800090c";
		wait for Clk_period;
		Addr <=  "00000110100111";
		Trees_din <= x"19008b08";
		wait for Clk_period;
		Addr <=  "00000110101000";
		Trees_din <= x"0000af04";
		wait for Clk_period;
		Addr <=  "00000110101001";
		Trees_din <= x"010a0765";
		wait for Clk_period;
		Addr <=  "00000110101010";
		Trees_din <= x"ffa20765";
		wait for Clk_period;
		Addr <=  "00000110101011";
		Trees_din <= x"ff880765";
		wait for Clk_period;
		Addr <=  "00000110101100";
		Trees_din <= x"1005e408";
		wait for Clk_period;
		Addr <=  "00000110101101";
		Trees_din <= x"1b002d04";
		wait for Clk_period;
		Addr <=  "00000110101110";
		Trees_din <= x"ffd30765";
		wait for Clk_period;
		Addr <=  "00000110101111";
		Trees_din <= x"ff620765";
		wait for Clk_period;
		Addr <=  "00000110110000";
		Trees_din <= x"1c003604";
		wait for Clk_period;
		Addr <=  "00000110110001";
		Trees_din <= x"ff8b0765";
		wait for Clk_period;
		Addr <=  "00000110110010";
		Trees_din <= x"005c0765";
		wait for Clk_period;
		Addr <=  "00000110110011";
		Trees_din <= x"06f50b04";
		wait for Clk_period;
		Addr <=  "00000110110100";
		Trees_din <= x"ff940765";
		wait for Clk_period;
		Addr <=  "00000110110101";
		Trees_din <= x"00c90765";
		wait for Clk_period;
		Addr <=  "00000110110110";
		Trees_din <= x"0307f524";
		wait for Clk_period;
		Addr <=  "00000110110111";
		Trees_din <= x"00f9b904";
		wait for Clk_period;
		Addr <=  "00000110111000";
		Trees_din <= x"ff6b0765";
		wait for Clk_period;
		Addr <=  "00000110111001";
		Trees_din <= x"12fe8310";
		wait for Clk_period;
		Addr <=  "00000110111010";
		Trees_din <= x"16018d08";
		wait for Clk_period;
		Addr <=  "00000110111011";
		Trees_din <= x"16001e04";
		wait for Clk_period;
		Addr <=  "00000110111100";
		Trees_din <= x"fffa0765";
		wait for Clk_period;
		Addr <=  "00000110111101";
		Trees_din <= x"ff7f0765";
		wait for Clk_period;
		Addr <=  "00000110111110";
		Trees_din <= x"0f000404";
		wait for Clk_period;
		Addr <=  "00000110111111";
		Trees_din <= x"ffeb0765";
		wait for Clk_period;
		Addr <=  "00000111000000";
		Trees_din <= x"00e80765";
		wait for Clk_period;
		Addr <=  "00000111000001";
		Trees_din <= x"0a028208";
		wait for Clk_period;
		Addr <=  "00000111000010";
		Trees_din <= x"05f92804";
		wait for Clk_period;
		Addr <=  "00000111000011";
		Trees_din <= x"ff910765";
		wait for Clk_period;
		Addr <=  "00000111000100";
		Trees_din <= x"00340765";
		wait for Clk_period;
		Addr <=  "00000111000101";
		Trees_din <= x"18004604";
		wait for Clk_period;
		Addr <=  "00000111000110";
		Trees_din <= x"ff7c0765";
		wait for Clk_period;
		Addr <=  "00000111000111";
		Trees_din <= x"00350765";
		wait for Clk_period;
		Addr <=  "00000111001000";
		Trees_din <= x"030fb414";
		wait for Clk_period;
		Addr <=  "00000111001001";
		Trees_din <= x"1500b110";
		wait for Clk_period;
		Addr <=  "00000111001010";
		Trees_din <= x"04041b08";
		wait for Clk_period;
		Addr <=  "00000111001011";
		Trees_din <= x"1702dc04";
		wait for Clk_period;
		Addr <=  "00000111001100";
		Trees_din <= x"00ae0765";
		wait for Clk_period;
		Addr <=  "00000111001101";
		Trees_din <= x"00300765";
		wait for Clk_period;
		Addr <=  "00000111001110";
		Trees_din <= x"08003504";
		wait for Clk_period;
		Addr <=  "00000111001111";
		Trees_din <= x"ffc30765";
		wait for Clk_period;
		Addr <=  "00000111010000";
		Trees_din <= x"00650765";
		wait for Clk_period;
		Addr <=  "00000111010001";
		Trees_din <= x"ff9d0765";
		wait for Clk_period;
		Addr <=  "00000111010010";
		Trees_din <= x"05f54504";
		wait for Clk_period;
		Addr <=  "00000111010011";
		Trees_din <= x"00450765";
		wait for Clk_period;
		Addr <=  "00000111010100";
		Trees_din <= x"08000a08";
		wait for Clk_period;
		Addr <=  "00000111010101";
		Trees_din <= x"0b046c04";
		wait for Clk_period;
		Addr <=  "00000111010110";
		Trees_din <= x"00980765";
		wait for Clk_period;
		Addr <=  "00000111010111";
		Trees_din <= x"ffc80765";
		wait for Clk_period;
		Addr <=  "00000111011000";
		Trees_din <= x"00c10765";
		wait for Clk_period;
		Addr <=  "00000111011001";
		Trees_din <= x"03029128";
		wait for Clk_period;
		Addr <=  "00000111011010";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00000111011011";
		Trees_din <= x"ff630841";
		wait for Clk_period;
		Addr <=  "00000111011100";
		Trees_din <= x"07005e1c";
		wait for Clk_period;
		Addr <=  "00000111011101";
		Trees_din <= x"0800090c";
		wait for Clk_period;
		Addr <=  "00000111011110";
		Trees_din <= x"19008b08";
		wait for Clk_period;
		Addr <=  "00000111011111";
		Trees_din <= x"0000af04";
		wait for Clk_period;
		Addr <=  "00000111100000";
		Trees_din <= x"00dd0841";
		wait for Clk_period;
		Addr <=  "00000111100001";
		Trees_din <= x"ffa70841";
		wait for Clk_period;
		Addr <=  "00000111100010";
		Trees_din <= x"ff8e0841";
		wait for Clk_period;
		Addr <=  "00000111100011";
		Trees_din <= x"0a041608";
		wait for Clk_period;
		Addr <=  "00000111100100";
		Trees_din <= x"03fe8b04";
		wait for Clk_period;
		Addr <=  "00000111100101";
		Trees_din <= x"00030841";
		wait for Clk_period;
		Addr <=  "00000111100110";
		Trees_din <= x"ff6c0841";
		wait for Clk_period;
		Addr <=  "00000111100111";
		Trees_din <= x"0a046704";
		wait for Clk_period;
		Addr <=  "00000111101000";
		Trees_din <= x"00a60841";
		wait for Clk_period;
		Addr <=  "00000111101001";
		Trees_din <= x"ff870841";
		wait for Clk_period;
		Addr <=  "00000111101010";
		Trees_din <= x"0efebe04";
		wait for Clk_period;
		Addr <=  "00000111101011";
		Trees_din <= x"00b90841";
		wait for Clk_period;
		Addr <=  "00000111101100";
		Trees_din <= x"ff990841";
		wait for Clk_period;
		Addr <=  "00000111101101";
		Trees_din <= x"0308a91c";
		wait for Clk_period;
		Addr <=  "00000111101110";
		Trees_din <= x"05f86604";
		wait for Clk_period;
		Addr <=  "00000111101111";
		Trees_din <= x"ff6d0841";
		wait for Clk_period;
		Addr <=  "00000111110000";
		Trees_din <= x"0101fc0c";
		wait for Clk_period;
		Addr <=  "00000111110001";
		Trees_din <= x"0203f908";
		wait for Clk_period;
		Addr <=  "00000111110010";
		Trees_din <= x"00fd2504";
		wait for Clk_period;
		Addr <=  "00000111110011";
		Trees_din <= x"ffb50841";
		wait for Clk_period;
		Addr <=  "00000111110100";
		Trees_din <= x"00310841";
		wait for Clk_period;
		Addr <=  "00000111110101";
		Trees_din <= x"ff6c0841";
		wait for Clk_period;
		Addr <=  "00000111110110";
		Trees_din <= x"1b004808";
		wait for Clk_period;
		Addr <=  "00000111110111";
		Trees_din <= x"06f5af04";
		wait for Clk_period;
		Addr <=  "00000111111000";
		Trees_din <= x"00860841";
		wait for Clk_period;
		Addr <=  "00000111111001";
		Trees_din <= x"ffe20841";
		wait for Clk_period;
		Addr <=  "00000111111010";
		Trees_din <= x"00f40841";
		wait for Clk_period;
		Addr <=  "00000111111011";
		Trees_din <= x"030fb41c";
		wait for Clk_period;
		Addr <=  "00000111111100";
		Trees_din <= x"06f5d010";
		wait for Clk_period;
		Addr <=  "00000111111101";
		Trees_din <= x"0d012208";
		wait for Clk_period;
		Addr <=  "00000111111110";
		Trees_din <= x"0d000704";
		wait for Clk_period;
		Addr <=  "00000111111111";
		Trees_din <= x"ffb90841";
		wait for Clk_period;
		Addr <=  "00001000000000";
		Trees_din <= x"00c10841";
		wait for Clk_period;
		Addr <=  "00001000000001";
		Trees_din <= x"1600e204";
		wait for Clk_period;
		Addr <=  "00001000000010";
		Trees_din <= x"008e0841";
		wait for Clk_period;
		Addr <=  "00001000000011";
		Trees_din <= x"ffc80841";
		wait for Clk_period;
		Addr <=  "00001000000100";
		Trees_din <= x"1500af08";
		wait for Clk_period;
		Addr <=  "00001000000101";
		Trees_din <= x"01fb7504";
		wait for Clk_period;
		Addr <=  "00001000000110";
		Trees_din <= x"00400841";
		wait for Clk_period;
		Addr <=  "00001000000111";
		Trees_din <= x"00a00841";
		wait for Clk_period;
		Addr <=  "00001000001000";
		Trees_din <= x"ffb40841";
		wait for Clk_period;
		Addr <=  "00001000001001";
		Trees_din <= x"05f54504";
		wait for Clk_period;
		Addr <=  "00001000001010";
		Trees_din <= x"00370841";
		wait for Clk_period;
		Addr <=  "00001000001011";
		Trees_din <= x"08000a08";
		wait for Clk_period;
		Addr <=  "00001000001100";
		Trees_din <= x"04065f04";
		wait for Clk_period;
		Addr <=  "00001000001101";
		Trees_din <= x"008a0841";
		wait for Clk_period;
		Addr <=  "00001000001110";
		Trees_din <= x"ffc80841";
		wait for Clk_period;
		Addr <=  "00001000001111";
		Trees_din <= x"00b50841";
		wait for Clk_period;
		Addr <=  "00001000010000";
		Trees_din <= x"03029128";
		wait for Clk_period;
		Addr <=  "00001000010001";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00001000010010";
		Trees_din <= x"ff64093d";
		wait for Clk_period;
		Addr <=  "00001000010011";
		Trees_din <= x"08000910";
		wait for Clk_period;
		Addr <=  "00001000010100";
		Trees_din <= x"08000508";
		wait for Clk_period;
		Addr <=  "00001000010101";
		Trees_din <= x"1603ed04";
		wait for Clk_period;
		Addr <=  "00001000010110";
		Trees_din <= x"ff8f093d";
		wait for Clk_period;
		Addr <=  "00001000010111";
		Trees_din <= x"0017093d";
		wait for Clk_period;
		Addr <=  "00001000011000";
		Trees_din <= x"0afc6404";
		wait for Clk_period;
		Addr <=  "00001000011001";
		Trees_din <= x"002e093d";
		wait for Clk_period;
		Addr <=  "00001000011010";
		Trees_din <= x"00c9093d";
		wait for Clk_period;
		Addr <=  "00001000011011";
		Trees_din <= x"07005e10";
		wait for Clk_period;
		Addr <=  "00001000011100";
		Trees_din <= x"1005e408";
		wait for Clk_period;
		Addr <=  "00001000011101";
		Trees_din <= x"1b002d04";
		wait for Clk_period;
		Addr <=  "00001000011110";
		Trees_din <= x"ffeb093d";
		wait for Clk_period;
		Addr <=  "00001000011111";
		Trees_din <= x"ff66093d";
		wait for Clk_period;
		Addr <=  "00001000100000";
		Trees_din <= x"0301b004";
		wait for Clk_period;
		Addr <=  "00001000100001";
		Trees_din <= x"ff98093d";
		wait for Clk_period;
		Addr <=  "00001000100010";
		Trees_din <= x"005f093d";
		wait for Clk_period;
		Addr <=  "00001000100011";
		Trees_din <= x"0034093d";
		wait for Clk_period;
		Addr <=  "00001000100100";
		Trees_din <= x"030bbf2c";
		wait for Clk_period;
		Addr <=  "00001000100101";
		Trees_din <= x"02053820";
		wait for Clk_period;
		Addr <=  "00001000100110";
		Trees_din <= x"15008210";
		wait for Clk_period;
		Addr <=  "00001000100111";
		Trees_din <= x"0bf9a008";
		wait for Clk_period;
		Addr <=  "00001000101000";
		Trees_din <= x"01036504";
		wait for Clk_period;
		Addr <=  "00001000101001";
		Trees_din <= x"000f093d";
		wait for Clk_period;
		Addr <=  "00001000101010";
		Trees_din <= x"00ab093d";
		wait for Clk_period;
		Addr <=  "00001000101011";
		Trees_din <= x"08011404";
		wait for Clk_period;
		Addr <=  "00001000101100";
		Trees_din <= x"ff5f093d";
		wait for Clk_period;
		Addr <=  "00001000101101";
		Trees_din <= x"0014093d";
		wait for Clk_period;
		Addr <=  "00001000101110";
		Trees_din <= x"03063408";
		wait for Clk_period;
		Addr <=  "00001000101111";
		Trees_din <= x"10fa2804";
		wait for Clk_period;
		Addr <=  "00001000110000";
		Trees_din <= x"ff74093d";
		wait for Clk_period;
		Addr <=  "00001000110001";
		Trees_din <= x"001b093d";
		wait for Clk_period;
		Addr <=  "00001000110010";
		Trees_din <= x"0400f004";
		wait for Clk_period;
		Addr <=  "00001000110011";
		Trees_din <= x"0089093d";
		wait for Clk_period;
		Addr <=  "00001000110100";
		Trees_din <= x"002c093d";
		wait for Clk_period;
		Addr <=  "00001000110101";
		Trees_din <= x"01037504";
		wait for Clk_period;
		Addr <=  "00001000110110";
		Trees_din <= x"ff6f093d";
		wait for Clk_period;
		Addr <=  "00001000110111";
		Trees_din <= x"0800bc04";
		wait for Clk_period;
		Addr <=  "00001000111000";
		Trees_din <= x"009f093d";
		wait for Clk_period;
		Addr <=  "00001000111001";
		Trees_din <= x"ffdc093d";
		wait for Clk_period;
		Addr <=  "00001000111010";
		Trees_din <= x"14004b14";
		wait for Clk_period;
		Addr <=  "00001000111011";
		Trees_din <= x"030fb40c";
		wait for Clk_period;
		Addr <=  "00001000111100";
		Trees_din <= x"17036004";
		wait for Clk_period;
		Addr <=  "00001000111101";
		Trees_din <= x"ff48093d";
		wait for Clk_period;
		Addr <=  "00001000111110";
		Trees_din <= x"06f7a804";
		wait for Clk_period;
		Addr <=  "00001000111111";
		Trees_din <= x"007e093d";
		wait for Clk_period;
		Addr <=  "00001001000000";
		Trees_din <= x"ffd7093d";
		wait for Clk_period;
		Addr <=  "00001001000001";
		Trees_din <= x"09005604";
		wait for Clk_period;
		Addr <=  "00001001000010";
		Trees_din <= x"0098093d";
		wait for Clk_period;
		Addr <=  "00001001000011";
		Trees_din <= x"0001093d";
		wait for Clk_period;
		Addr <=  "00001001000100";
		Trees_din <= x"1104d510";
		wait for Clk_period;
		Addr <=  "00001001000101";
		Trees_din <= x"1900a608";
		wait for Clk_period;
		Addr <=  "00001001000110";
		Trees_din <= x"0c03bc04";
		wait for Clk_period;
		Addr <=  "00001001000111";
		Trees_din <= x"00b0093d";
		wait for Clk_period;
		Addr <=  "00001001001000";
		Trees_din <= x"0001093d";
		wait for Clk_period;
		Addr <=  "00001001001001";
		Trees_din <= x"1e005e04";
		wait for Clk_period;
		Addr <=  "00001001001010";
		Trees_din <= x"007e093d";
		wait for Clk_period;
		Addr <=  "00001001001011";
		Trees_din <= x"ff6c093d";
		wait for Clk_period;
		Addr <=  "00001001001100";
		Trees_din <= x"00fae404";
		wait for Clk_period;
		Addr <=  "00001001001101";
		Trees_din <= x"ff92093d";
		wait for Clk_period;
		Addr <=  "00001001001110";
		Trees_din <= x"0074093d";
		wait for Clk_period;
		Addr <=  "00001001001111";
		Trees_din <= x"0302912c";
		wait for Clk_period;
		Addr <=  "00001001010000";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00001001010001";
		Trees_din <= x"ff650a49";
		wait for Clk_period;
		Addr <=  "00001001010010";
		Trees_din <= x"08007118";
		wait for Clk_period;
		Addr <=  "00001001010011";
		Trees_din <= x"11000d0c";
		wait for Clk_period;
		Addr <=  "00001001010100";
		Trees_din <= x"06f59704";
		wait for Clk_period;
		Addr <=  "00001001010101";
		Trees_din <= x"ff9d0a49";
		wait for Clk_period;
		Addr <=  "00001001010110";
		Trees_din <= x"02016004";
		wait for Clk_period;
		Addr <=  "00001001010111";
		Trees_din <= x"000b0a49";
		wait for Clk_period;
		Addr <=  "00001001011000";
		Trees_din <= x"01310a49";
		wait for Clk_period;
		Addr <=  "00001001011001";
		Trees_din <= x"1a00b008";
		wait for Clk_period;
		Addr <=  "00001001011010";
		Trees_din <= x"0000af04";
		wait for Clk_period;
		Addr <=  "00001001011011";
		Trees_din <= x"00800a49";
		wait for Clk_period;
		Addr <=  "00001001011100";
		Trees_din <= x"ff9b0a49";
		wait for Clk_period;
		Addr <=  "00001001011101";
		Trees_din <= x"ff780a49";
		wait for Clk_period;
		Addr <=  "00001001011110";
		Trees_din <= x"0a041608";
		wait for Clk_period;
		Addr <=  "00001001011111";
		Trees_din <= x"0ef94304";
		wait for Clk_period;
		Addr <=  "00001001100000";
		Trees_din <= x"000c0a49";
		wait for Clk_period;
		Addr <=  "00001001100001";
		Trees_din <= x"ff680a49";
		wait for Clk_period;
		Addr <=  "00001001100010";
		Trees_din <= x"0a046704";
		wait for Clk_period;
		Addr <=  "00001001100011";
		Trees_din <= x"00ab0a49";
		wait for Clk_period;
		Addr <=  "00001001100100";
		Trees_din <= x"ff930a49";
		wait for Clk_period;
		Addr <=  "00001001100101";
		Trees_din <= x"030bbf34";
		wait for Clk_period;
		Addr <=  "00001001100110";
		Trees_din <= x"09004e20";
		wait for Clk_period;
		Addr <=  "00001001100111";
		Trees_din <= x"0d011510";
		wait for Clk_period;
		Addr <=  "00001001101000";
		Trees_din <= x"0f003708";
		wait for Clk_period;
		Addr <=  "00001001101001";
		Trees_din <= x"1b003104";
		wait for Clk_period;
		Addr <=  "00001001101010";
		Trees_din <= x"00530a49";
		wait for Clk_period;
		Addr <=  "00001001101011";
		Trees_din <= x"00fb0a49";
		wait for Clk_period;
		Addr <=  "00001001101100";
		Trees_din <= x"0c00a004";
		wait for Clk_period;
		Addr <=  "00001001101101";
		Trees_din <= x"ffbf0a49";
		wait for Clk_period;
		Addr <=  "00001001101110";
		Trees_din <= x"007b0a49";
		wait for Clk_period;
		Addr <=  "00001001101111";
		Trees_din <= x"0405b608";
		wait for Clk_period;
		Addr <=  "00001001110000";
		Trees_din <= x"1d003e04";
		wait for Clk_period;
		Addr <=  "00001001110001";
		Trees_din <= x"ff8c0a49";
		wait for Clk_period;
		Addr <=  "00001001110010";
		Trees_din <= x"00380a49";
		wait for Clk_period;
		Addr <=  "00001001110011";
		Trees_din <= x"10facc04";
		wait for Clk_period;
		Addr <=  "00001001110100";
		Trees_din <= x"00b00a49";
		wait for Clk_period;
		Addr <=  "00001001110101";
		Trees_din <= x"00140a49";
		wait for Clk_period;
		Addr <=  "00001001110110";
		Trees_din <= x"0c002904";
		wait for Clk_period;
		Addr <=  "00001001110111";
		Trees_din <= x"ff660a49";
		wait for Clk_period;
		Addr <=  "00001001111000";
		Trees_din <= x"09005208";
		wait for Clk_period;
		Addr <=  "00001001111001";
		Trees_din <= x"1500a404";
		wait for Clk_period;
		Addr <=  "00001001111010";
		Trees_din <= x"ff8d0a49";
		wait for Clk_period;
		Addr <=  "00001001111011";
		Trees_din <= x"00190a49";
		wait for Clk_period;
		Addr <=  "00001001111100";
		Trees_din <= x"0101c604";
		wait for Clk_period;
		Addr <=  "00001001111101";
		Trees_din <= x"00080a49";
		wait for Clk_period;
		Addr <=  "00001001111110";
		Trees_din <= x"005a0a49";
		wait for Clk_period;
		Addr <=  "00001001111111";
		Trees_din <= x"14004b10";
		wait for Clk_period;
		Addr <=  "00001010000000";
		Trees_din <= x"01f9cb04";
		wait for Clk_period;
		Addr <=  "00001010000001";
		Trees_din <= x"00900a49";
		wait for Clk_period;
		Addr <=  "00001010000010";
		Trees_din <= x"04fe3404";
		wait for Clk_period;
		Addr <=  "00001010000011";
		Trees_din <= x"ff690a49";
		wait for Clk_period;
		Addr <=  "00001010000100";
		Trees_din <= x"0404aa04";
		wait for Clk_period;
		Addr <=  "00001010000101";
		Trees_din <= x"00820a49";
		wait for Clk_period;
		Addr <=  "00001010000110";
		Trees_din <= x"ff920a49";
		wait for Clk_period;
		Addr <=  "00001010000111";
		Trees_din <= x"0407e10c";
		wait for Clk_period;
		Addr <=  "00001010001000";
		Trees_din <= x"18003708";
		wait for Clk_period;
		Addr <=  "00001010001001";
		Trees_din <= x"18003704";
		wait for Clk_period;
		Addr <=  "00001010001010";
		Trees_din <= x"00900a49";
		wait for Clk_period;
		Addr <=  "00001010001011";
		Trees_din <= x"ff890a49";
		wait for Clk_period;
		Addr <=  "00001010001100";
		Trees_din <= x"00ac0a49";
		wait for Clk_period;
		Addr <=  "00001010001101";
		Trees_din <= x"0c03bc08";
		wait for Clk_period;
		Addr <=  "00001010001110";
		Trees_din <= x"02001704";
		wait for Clk_period;
		Addr <=  "00001010001111";
		Trees_din <= x"008b0a49";
		wait for Clk_period;
		Addr <=  "00001010010000";
		Trees_din <= x"ffdd0a49";
		wait for Clk_period;
		Addr <=  "00001010010001";
		Trees_din <= x"ffa60a49";
		wait for Clk_period;
		Addr <=  "00001010010010";
		Trees_din <= x"0301f920";
		wait for Clk_period;
		Addr <=  "00001010010011";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00001010010100";
		Trees_din <= x"ff650b25";
		wait for Clk_period;
		Addr <=  "00001010010101";
		Trees_din <= x"07005e14";
		wait for Clk_period;
		Addr <=  "00001010010110";
		Trees_din <= x"0d03ab0c";
		wait for Clk_period;
		Addr <=  "00001010010111";
		Trees_din <= x"11036904";
		wait for Clk_period;
		Addr <=  "00001010011000";
		Trees_din <= x"ff6a0b25";
		wait for Clk_period;
		Addr <=  "00001010011001";
		Trees_din <= x"0bfad604";
		wait for Clk_period;
		Addr <=  "00001010011010";
		Trees_din <= x"009e0b25";
		wait for Clk_period;
		Addr <=  "00001010011011";
		Trees_din <= x"ff920b25";
		wait for Clk_period;
		Addr <=  "00001010011100";
		Trees_din <= x"1700b204";
		wait for Clk_period;
		Addr <=  "00001010011101";
		Trees_din <= x"ff9f0b25";
		wait for Clk_period;
		Addr <=  "00001010011110";
		Trees_din <= x"00b50b25";
		wait for Clk_period;
		Addr <=  "00001010011111";
		Trees_din <= x"0202b804";
		wait for Clk_period;
		Addr <=  "00001010100000";
		Trees_din <= x"ffa50b25";
		wait for Clk_period;
		Addr <=  "00001010100001";
		Trees_din <= x"009a0b25";
		wait for Clk_period;
		Addr <=  "00001010100010";
		Trees_din <= x"0308a924";
		wait for Clk_period;
		Addr <=  "00001010100011";
		Trees_din <= x"05f86604";
		wait for Clk_period;
		Addr <=  "00001010100100";
		Trees_din <= x"ff730b25";
		wait for Clk_period;
		Addr <=  "00001010100101";
		Trees_din <= x"0c01c810";
		wait for Clk_period;
		Addr <=  "00001010100110";
		Trees_din <= x"0101d108";
		wait for Clk_period;
		Addr <=  "00001010100111";
		Trees_din <= x"00001404";
		wait for Clk_period;
		Addr <=  "00001010101000";
		Trees_din <= x"ffc80b25";
		wait for Clk_period;
		Addr <=  "00001010101001";
		Trees_din <= x"003e0b25";
		wait for Clk_period;
		Addr <=  "00001010101010";
		Trees_din <= x"11028004";
		wait for Clk_period;
		Addr <=  "00001010101011";
		Trees_din <= x"009e0b25";
		wait for Clk_period;
		Addr <=  "00001010101100";
		Trees_din <= x"fff70b25";
		wait for Clk_period;
		Addr <=  "00001010101101";
		Trees_din <= x"0f012e08";
		wait for Clk_period;
		Addr <=  "00001010101110";
		Trees_din <= x"09005804";
		wait for Clk_period;
		Addr <=  "00001010101111";
		Trees_din <= x"002c0b25";
		wait for Clk_period;
		Addr <=  "00001010110000";
		Trees_din <= x"ff990b25";
		wait for Clk_period;
		Addr <=  "00001010110001";
		Trees_din <= x"13ffc104";
		wait for Clk_period;
		Addr <=  "00001010110010";
		Trees_din <= x"ffdb0b25";
		wait for Clk_period;
		Addr <=  "00001010110011";
		Trees_din <= x"ff5e0b25";
		wait for Clk_period;
		Addr <=  "00001010110100";
		Trees_din <= x"030fb420";
		wait for Clk_period;
		Addr <=  "00001010110101";
		Trees_din <= x"01fdeb10";
		wait for Clk_period;
		Addr <=  "00001010110110";
		Trees_din <= x"01fd0908";
		wait for Clk_period;
		Addr <=  "00001010110111";
		Trees_din <= x"1a00a104";
		wait for Clk_period;
		Addr <=  "00001010111000";
		Trees_din <= x"ff930b25";
		wait for Clk_period;
		Addr <=  "00001010111001";
		Trees_din <= x"00550b25";
		wait for Clk_period;
		Addr <=  "00001010111010";
		Trees_din <= x"04041b04";
		wait for Clk_period;
		Addr <=  "00001010111011";
		Trees_din <= x"00250b25";
		wait for Clk_period;
		Addr <=  "00001010111100";
		Trees_din <= x"ff5c0b25";
		wait for Clk_period;
		Addr <=  "00001010111101";
		Trees_din <= x"0d029108";
		wait for Clk_period;
		Addr <=  "00001010111110";
		Trees_din <= x"00f8f604";
		wait for Clk_period;
		Addr <=  "00001010111111";
		Trees_din <= x"00320b25";
		wait for Clk_period;
		Addr <=  "00001011000000";
		Trees_din <= x"00bb0b25";
		wait for Clk_period;
		Addr <=  "00001011000001";
		Trees_din <= x"0d030704";
		wait for Clk_period;
		Addr <=  "00001011000010";
		Trees_din <= x"ff610b25";
		wait for Clk_period;
		Addr <=  "00001011000011";
		Trees_din <= x"00630b25";
		wait for Clk_period;
		Addr <=  "00001011000100";
		Trees_din <= x"08002508";
		wait for Clk_period;
		Addr <=  "00001011000101";
		Trees_din <= x"0f009a04";
		wait for Clk_period;
		Addr <=  "00001011000110";
		Trees_din <= x"ffac0b25";
		wait for Clk_period;
		Addr <=  "00001011000111";
		Trees_din <= x"00810b25";
		wait for Clk_period;
		Addr <=  "00001011001000";
		Trees_din <= x"00a20b25";
		wait for Clk_period;
		Addr <=  "00001011001001";
		Trees_din <= x"0301f920";
		wait for Clk_period;
		Addr <=  "00001011001010";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00001011001011";
		Trees_din <= x"ff660c01";
		wait for Clk_period;
		Addr <=  "00001011001100";
		Trees_din <= x"02031008";
		wait for Clk_period;
		Addr <=  "00001011001101";
		Trees_din <= x"0a041604";
		wait for Clk_period;
		Addr <=  "00001011001110";
		Trees_din <= x"ff6d0c01";
		wait for Clk_period;
		Addr <=  "00001011001111";
		Trees_din <= x"001c0c01";
		wait for Clk_period;
		Addr <=  "00001011010000";
		Trees_din <= x"0800710c";
		wait for Clk_period;
		Addr <=  "00001011010001";
		Trees_din <= x"05faba04";
		wait for Clk_period;
		Addr <=  "00001011010010";
		Trees_din <= x"ffa50c01";
		wait for Clk_period;
		Addr <=  "00001011010011";
		Trees_din <= x"01027d04";
		wait for Clk_period;
		Addr <=  "00001011010100";
		Trees_din <= x"fff80c01";
		wait for Clk_period;
		Addr <=  "00001011010101";
		Trees_din <= x"01010c01";
		wait for Clk_period;
		Addr <=  "00001011010110";
		Trees_din <= x"0d006b04";
		wait for Clk_period;
		Addr <=  "00001011010111";
		Trees_din <= x"00210c01";
		wait for Clk_period;
		Addr <=  "00001011011000";
		Trees_din <= x"ff800c01";
		wait for Clk_period;
		Addr <=  "00001011011001";
		Trees_din <= x"0308a924";
		wait for Clk_period;
		Addr <=  "00001011011010";
		Trees_din <= x"05f86604";
		wait for Clk_period;
		Addr <=  "00001011011011";
		Trees_din <= x"ff780c01";
		wait for Clk_period;
		Addr <=  "00001011011100";
		Trees_din <= x"0c01c810";
		wait for Clk_period;
		Addr <=  "00001011011101";
		Trees_din <= x"0101d108";
		wait for Clk_period;
		Addr <=  "00001011011110";
		Trees_din <= x"00001404";
		wait for Clk_period;
		Addr <=  "00001011011111";
		Trees_din <= x"ffcf0c01";
		wait for Clk_period;
		Addr <=  "00001011100000";
		Trees_din <= x"00340c01";
		wait for Clk_period;
		Addr <=  "00001011100001";
		Trees_din <= x"15009804";
		wait for Clk_period;
		Addr <=  "00001011100010";
		Trees_din <= x"008e0c01";
		wait for Clk_period;
		Addr <=  "00001011100011";
		Trees_din <= x"fffe0c01";
		wait for Clk_period;
		Addr <=  "00001011100100";
		Trees_din <= x"06f54908";
		wait for Clk_period;
		Addr <=  "00001011100101";
		Trees_din <= x"11fd4604";
		wait for Clk_period;
		Addr <=  "00001011100110";
		Trees_din <= x"001a0c01";
		wait for Clk_period;
		Addr <=  "00001011100111";
		Trees_din <= x"ff6b0c01";
		wait for Clk_period;
		Addr <=  "00001011101000";
		Trees_din <= x"0305c704";
		wait for Clk_period;
		Addr <=  "00001011101001";
		Trees_din <= x"ffcc0c01";
		wait for Clk_period;
		Addr <=  "00001011101010";
		Trees_din <= x"00340c01";
		wait for Clk_period;
		Addr <=  "00001011101011";
		Trees_din <= x"030fb420";
		wait for Clk_period;
		Addr <=  "00001011101100";
		Trees_din <= x"01fdeb10";
		wait for Clk_period;
		Addr <=  "00001011101101";
		Trees_din <= x"01fd0908";
		wait for Clk_period;
		Addr <=  "00001011101110";
		Trees_din <= x"1a00a104";
		wait for Clk_period;
		Addr <=  "00001011101111";
		Trees_din <= x"ffa10c01";
		wait for Clk_period;
		Addr <=  "00001011110000";
		Trees_din <= x"00490c01";
		wait for Clk_period;
		Addr <=  "00001011110001";
		Trees_din <= x"0d017e04";
		wait for Clk_period;
		Addr <=  "00001011110010";
		Trees_din <= x"00390c01";
		wait for Clk_period;
		Addr <=  "00001011110011";
		Trees_din <= x"ff710c01";
		wait for Clk_period;
		Addr <=  "00001011110100";
		Trees_din <= x"0d029108";
		wait for Clk_period;
		Addr <=  "00001011110101";
		Trees_din <= x"00f8f604";
		wait for Clk_period;
		Addr <=  "00001011110110";
		Trees_din <= x"002c0c01";
		wait for Clk_period;
		Addr <=  "00001011110111";
		Trees_din <= x"00b00c01";
		wait for Clk_period;
		Addr <=  "00001011111000";
		Trees_din <= x"16032804";
		wait for Clk_period;
		Addr <=  "00001011111001";
		Trees_din <= x"006c0c01";
		wait for Clk_period;
		Addr <=  "00001011111010";
		Trees_din <= x"ff870c01";
		wait for Clk_period;
		Addr <=  "00001011111011";
		Trees_din <= x"08002508";
		wait for Clk_period;
		Addr <=  "00001011111100";
		Trees_din <= x"0f009a04";
		wait for Clk_period;
		Addr <=  "00001011111101";
		Trees_din <= x"ffae0c01";
		wait for Clk_period;
		Addr <=  "00001011111110";
		Trees_din <= x"00790c01";
		wait for Clk_period;
		Addr <=  "00001011111111";
		Trees_din <= x"009d0c01";
		wait for Clk_period;
		Addr <=  "00001100000000";
		Trees_din <= x"0301f920";
		wait for Clk_period;
		Addr <=  "00001100000001";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00001100000010";
		Trees_din <= x"ff670cf5";
		wait for Clk_period;
		Addr <=  "00001100000011";
		Trees_din <= x"02031008";
		wait for Clk_period;
		Addr <=  "00001100000100";
		Trees_din <= x"05f89e04";
		wait for Clk_period;
		Addr <=  "00001100000101";
		Trees_din <= x"00240cf5";
		wait for Clk_period;
		Addr <=  "00001100000110";
		Trees_din <= x"ff6f0cf5";
		wait for Clk_period;
		Addr <=  "00001100000111";
		Trees_din <= x"0800710c";
		wait for Clk_period;
		Addr <=  "00001100001000";
		Trees_din <= x"05faba04";
		wait for Clk_period;
		Addr <=  "00001100001001";
		Trees_din <= x"ffaa0cf5";
		wait for Clk_period;
		Addr <=  "00001100001010";
		Trees_din <= x"01027d04";
		wait for Clk_period;
		Addr <=  "00001100001011";
		Trees_din <= x"fffa0cf5";
		wait for Clk_period;
		Addr <=  "00001100001100";
		Trees_din <= x"00da0cf5";
		wait for Clk_period;
		Addr <=  "00001100001101";
		Trees_din <= x"07005b04";
		wait for Clk_period;
		Addr <=  "00001100001110";
		Trees_din <= x"ff840cf5";
		wait for Clk_period;
		Addr <=  "00001100001111";
		Trees_din <= x"00240cf5";
		wait for Clk_period;
		Addr <=  "00001100010000";
		Trees_din <= x"030bbf38";
		wait for Clk_period;
		Addr <=  "00001100010001";
		Trees_din <= x"1100a21c";
		wait for Clk_period;
		Addr <=  "00001100010010";
		Trees_din <= x"1a00c910";
		wait for Clk_period;
		Addr <=  "00001100010011";
		Trees_din <= x"07005908";
		wait for Clk_period;
		Addr <=  "00001100010100";
		Trees_din <= x"09005a04";
		wait for Clk_period;
		Addr <=  "00001100010101";
		Trees_din <= x"ff700cf5";
		wait for Clk_period;
		Addr <=  "00001100010110";
		Trees_din <= x"00250cf5";
		wait for Clk_period;
		Addr <=  "00001100010111";
		Trees_din <= x"03063404";
		wait for Clk_period;
		Addr <=  "00001100011000";
		Trees_din <= x"fff00cf5";
		wait for Clk_period;
		Addr <=  "00001100011001";
		Trees_din <= x"008b0cf5";
		wait for Clk_period;
		Addr <=  "00001100011010";
		Trees_din <= x"0f000604";
		wait for Clk_period;
		Addr <=  "00001100011011";
		Trees_din <= x"ff770cf5";
		wait for Clk_period;
		Addr <=  "00001100011100";
		Trees_din <= x"11fdfc04";
		wait for Clk_period;
		Addr <=  "00001100011101";
		Trees_din <= x"fffb0cf5";
		wait for Clk_period;
		Addr <=  "00001100011110";
		Trees_din <= x"00a60cf5";
		wait for Clk_period;
		Addr <=  "00001100011111";
		Trees_din <= x"0303820c";
		wait for Clk_period;
		Addr <=  "00001100100000";
		Trees_din <= x"1603fe08";
		wait for Clk_period;
		Addr <=  "00001100100001";
		Trees_din <= x"1c002704";
		wait for Clk_period;
		Addr <=  "00001100100010";
		Trees_din <= x"001a0cf5";
		wait for Clk_period;
		Addr <=  "00001100100011";
		Trees_din <= x"ff680cf5";
		wait for Clk_period;
		Addr <=  "00001100100100";
		Trees_din <= x"00980cf5";
		wait for Clk_period;
		Addr <=  "00001100100101";
		Trees_din <= x"1a00c308";
		wait for Clk_period;
		Addr <=  "00001100100110";
		Trees_din <= x"0101a504";
		wait for Clk_period;
		Addr <=  "00001100100111";
		Trees_din <= x"00090cf5";
		wait for Clk_period;
		Addr <=  "00001100101000";
		Trees_din <= x"00b20cf5";
		wait for Clk_period;
		Addr <=  "00001100101001";
		Trees_din <= x"1e006704";
		wait for Clk_period;
		Addr <=  "00001100101010";
		Trees_din <= x"fffe0cf5";
		wait for Clk_period;
		Addr <=  "00001100101011";
		Trees_din <= x"ff7a0cf5";
		wait for Clk_period;
		Addr <=  "00001100101100";
		Trees_din <= x"14004b10";
		wait for Clk_period;
		Addr <=  "00001100101101";
		Trees_din <= x"01f9cb04";
		wait for Clk_period;
		Addr <=  "00001100101110";
		Trees_din <= x"007a0cf5";
		wait for Clk_period;
		Addr <=  "00001100101111";
		Trees_din <= x"04fe3404";
		wait for Clk_period;
		Addr <=  "00001100110000";
		Trees_din <= x"ff6f0cf5";
		wait for Clk_period;
		Addr <=  "00001100110001";
		Trees_din <= x"0404aa04";
		wait for Clk_period;
		Addr <=  "00001100110010";
		Trees_din <= x"006c0cf5";
		wait for Clk_period;
		Addr <=  "00001100110011";
		Trees_din <= x"ff9a0cf5";
		wait for Clk_period;
		Addr <=  "00001100110100";
		Trees_din <= x"1104d510";
		wait for Clk_period;
		Addr <=  "00001100110101";
		Trees_din <= x"1900a608";
		wait for Clk_period;
		Addr <=  "00001100110110";
		Trees_din <= x"0a077a04";
		wait for Clk_period;
		Addr <=  "00001100110111";
		Trees_din <= x"00990cf5";
		wait for Clk_period;
		Addr <=  "00001100111000";
		Trees_din <= x"ffe50cf5";
		wait for Clk_period;
		Addr <=  "00001100111001";
		Trees_din <= x"16033104";
		wait for Clk_period;
		Addr <=  "00001100111010";
		Trees_din <= x"00840cf5";
		wait for Clk_period;
		Addr <=  "00001100111011";
		Trees_din <= x"ffa50cf5";
		wait for Clk_period;
		Addr <=  "00001100111100";
		Trees_din <= x"ffdb0cf5";
		wait for Clk_period;
		Addr <=  "00001100111101";
		Trees_din <= x"0300490c";
		wait for Clk_period;
		Addr <=  "00001100111110";
		Trees_din <= x"00fcaf04";
		wait for Clk_period;
		Addr <=  "00001100111111";
		Trees_din <= x"00150db9";
		wait for Clk_period;
		Addr <=  "00001101000000";
		Trees_din <= x"1f005f04";
		wait for Clk_period;
		Addr <=  "00001101000001";
		Trees_din <= x"ff6a0db9";
		wait for Clk_period;
		Addr <=  "00001101000010";
		Trees_din <= x"00180db9";
		wait for Clk_period;
		Addr <=  "00001101000011";
		Trees_din <= x"0308a928";
		wait for Clk_period;
		Addr <=  "00001101000100";
		Trees_din <= x"18003308";
		wait for Clk_period;
		Addr <=  "00001101000101";
		Trees_din <= x"0b043104";
		wait for Clk_period;
		Addr <=  "00001101000110";
		Trees_din <= x"ff680db9";
		wait for Clk_period;
		Addr <=  "00001101000111";
		Trees_din <= x"00160db9";
		wait for Clk_period;
		Addr <=  "00001101001000";
		Trees_din <= x"1900a910";
		wait for Clk_period;
		Addr <=  "00001101001001";
		Trees_din <= x"00fd6408";
		wait for Clk_period;
		Addr <=  "00001101001010";
		Trees_din <= x"1a00b204";
		wait for Clk_period;
		Addr <=  "00001101001011";
		Trees_din <= x"00080db9";
		wait for Clk_period;
		Addr <=  "00001101001100";
		Trees_din <= x"ff8b0db9";
		wait for Clk_period;
		Addr <=  "00001101001101";
		Trees_din <= x"07005604";
		wait for Clk_period;
		Addr <=  "00001101001110";
		Trees_din <= x"ffc60db9";
		wait for Clk_period;
		Addr <=  "00001101001111";
		Trees_din <= x"00270db9";
		wait for Clk_period;
		Addr <=  "00001101010000";
		Trees_din <= x"1900b308";
		wait for Clk_period;
		Addr <=  "00001101010001";
		Trees_din <= x"07005604";
		wait for Clk_period;
		Addr <=  "00001101010010";
		Trees_din <= x"00bf0db9";
		wait for Clk_period;
		Addr <=  "00001101010011";
		Trees_din <= x"000d0db9";
		wait for Clk_period;
		Addr <=  "00001101010100";
		Trees_din <= x"10027a04";
		wait for Clk_period;
		Addr <=  "00001101010101";
		Trees_din <= x"00230db9";
		wait for Clk_period;
		Addr <=  "00001101010110";
		Trees_din <= x"ff840db9";
		wait for Clk_period;
		Addr <=  "00001101010111";
		Trees_din <= x"09004f10";
		wait for Clk_period;
		Addr <=  "00001101011000";
		Trees_din <= x"1500b10c";
		wait for Clk_period;
		Addr <=  "00001101011001";
		Trees_din <= x"14002d04";
		wait for Clk_period;
		Addr <=  "00001101011010";
		Trees_din <= x"fff00db9";
		wait for Clk_period;
		Addr <=  "00001101011011";
		Trees_din <= x"01006f04";
		wait for Clk_period;
		Addr <=  "00001101011100";
		Trees_din <= x"00a90db9";
		wait for Clk_period;
		Addr <=  "00001101011101";
		Trees_din <= x"00120db9";
		wait for Clk_period;
		Addr <=  "00001101011110";
		Trees_din <= x"ffed0db9";
		wait for Clk_period;
		Addr <=  "00001101011111";
		Trees_din <= x"04032b10";
		wait for Clk_period;
		Addr <=  "00001101100000";
		Trees_din <= x"09005008";
		wait for Clk_period;
		Addr <=  "00001101100001";
		Trees_din <= x"1e006904";
		wait for Clk_period;
		Addr <=  "00001101100010";
		Trees_din <= x"001e0db9";
		wait for Clk_period;
		Addr <=  "00001101100011";
		Trees_din <= x"ff820db9";
		wait for Clk_period;
		Addr <=  "00001101100100";
		Trees_din <= x"14004304";
		wait for Clk_period;
		Addr <=  "00001101100101";
		Trees_din <= x"000a0db9";
		wait for Clk_period;
		Addr <=  "00001101100110";
		Trees_din <= x"008f0db9";
		wait for Clk_period;
		Addr <=  "00001101100111";
		Trees_din <= x"02fe8308";
		wait for Clk_period;
		Addr <=  "00001101101000";
		Trees_din <= x"1d005404";
		wait for Clk_period;
		Addr <=  "00001101101001";
		Trees_din <= x"004c0db9";
		wait for Clk_period;
		Addr <=  "00001101101010";
		Trees_din <= x"ffbc0db9";
		wait for Clk_period;
		Addr <=  "00001101101011";
		Trees_din <= x"00fe2904";
		wait for Clk_period;
		Addr <=  "00001101101100";
		Trees_din <= x"00020db9";
		wait for Clk_period;
		Addr <=  "00001101101101";
		Trees_din <= x"ff600db9";
		wait for Clk_period;
		Addr <=  "00001101101110";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00001101101111";
		Trees_din <= x"03004914";
		wait for Clk_period;
		Addr <=  "00001101110000";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00001101110001";
		Trees_din <= x"ff680e89";
		wait for Clk_period;
		Addr <=  "00001101110010";
		Trees_din <= x"0800550c";
		wait for Clk_period;
		Addr <=  "00001101110011";
		Trees_din <= x"02031004";
		wait for Clk_period;
		Addr <=  "00001101110100";
		Trees_din <= x"ffa50e89";
		wait for Clk_period;
		Addr <=  "00001101110101";
		Trees_din <= x"07005804";
		wait for Clk_period;
		Addr <=  "00001101110110";
		Trees_din <= x"00c70e89";
		wait for Clk_period;
		Addr <=  "00001101110111";
		Trees_din <= x"00030e89";
		wait for Clk_period;
		Addr <=  "00001101111000";
		Trees_din <= x"ff7d0e89";
		wait for Clk_period;
		Addr <=  "00001101111001";
		Trees_din <= x"030bbf30";
		wait for Clk_period;
		Addr <=  "00001101111010";
		Trees_din <= x"02053820";
		wait for Clk_period;
		Addr <=  "00001101111011";
		Trees_din <= x"15008c10";
		wait for Clk_period;
		Addr <=  "00001101111100";
		Trees_din <= x"06f5d008";
		wait for Clk_period;
		Addr <=  "00001101111101";
		Trees_din <= x"06f37104";
		wait for Clk_period;
		Addr <=  "00001101111110";
		Trees_din <= x"002e0e89";
		wait for Clk_period;
		Addr <=  "00001101111111";
		Trees_din <= x"ff570e89";
		wait for Clk_period;
		Addr <=  "00001110000000";
		Trees_din <= x"11013d04";
		wait for Clk_period;
		Addr <=  "00001110000001";
		Trees_din <= x"ffaf0e89";
		wait for Clk_period;
		Addr <=  "00001110000010";
		Trees_din <= x"00360e89";
		wait for Clk_period;
		Addr <=  "00001110000011";
		Trees_din <= x"1100f508";
		wait for Clk_period;
		Addr <=  "00001110000100";
		Trees_din <= x"0f000404";
		wait for Clk_period;
		Addr <=  "00001110000101";
		Trees_din <= x"ff8f0e89";
		wait for Clk_period;
		Addr <=  "00001110000110";
		Trees_din <= x"00570e89";
		wait for Clk_period;
		Addr <=  "00001110000111";
		Trees_din <= x"18004204";
		wait for Clk_period;
		Addr <=  "00001110001000";
		Trees_din <= x"ffe10e89";
		wait for Clk_period;
		Addr <=  "00001110001001";
		Trees_din <= x"00430e89";
		wait for Clk_period;
		Addr <=  "00001110001010";
		Trees_din <= x"15008908";
		wait for Clk_period;
		Addr <=  "00001110001011";
		Trees_din <= x"14002004";
		wait for Clk_period;
		Addr <=  "00001110001100";
		Trees_din <= x"00760e89";
		wait for Clk_period;
		Addr <=  "00001110001101";
		Trees_din <= x"ffda0e89";
		wait for Clk_period;
		Addr <=  "00001110001110";
		Trees_din <= x"10f99904";
		wait for Clk_period;
		Addr <=  "00001110001111";
		Trees_din <= x"fff00e89";
		wait for Clk_period;
		Addr <=  "00001110010000";
		Trees_din <= x"ff730e89";
		wait for Clk_period;
		Addr <=  "00001110010001";
		Trees_din <= x"19009b10";
		wait for Clk_period;
		Addr <=  "00001110010010";
		Trees_din <= x"05f54504";
		wait for Clk_period;
		Addr <=  "00001110010011";
		Trees_din <= x"ffb70e89";
		wait for Clk_period;
		Addr <=  "00001110010100";
		Trees_din <= x"15007504";
		wait for Clk_period;
		Addr <=  "00001110010101";
		Trees_din <= x"ffde0e89";
		wait for Clk_period;
		Addr <=  "00001110010110";
		Trees_din <= x"0e041104";
		wait for Clk_period;
		Addr <=  "00001110010111";
		Trees_din <= x"00900e89";
		wait for Clk_period;
		Addr <=  "00001110011000";
		Trees_din <= x"fff40e89";
		wait for Clk_period;
		Addr <=  "00001110011001";
		Trees_din <= x"16033108";
		wait for Clk_period;
		Addr <=  "00001110011010";
		Trees_din <= x"0afc7c04";
		wait for Clk_period;
		Addr <=  "00001110011011";
		Trees_din <= x"fff10e89";
		wait for Clk_period;
		Addr <=  "00001110011100";
		Trees_din <= x"00860e89";
		wait for Clk_period;
		Addr <=  "00001110011101";
		Trees_din <= x"12028508";
		wait for Clk_period;
		Addr <=  "00001110011110";
		Trees_din <= x"0c00c704";
		wait for Clk_period;
		Addr <=  "00001110011111";
		Trees_din <= x"00180e89";
		wait for Clk_period;
		Addr <=  "00001110100000";
		Trees_din <= x"ff790e89";
		wait for Clk_period;
		Addr <=  "00001110100001";
		Trees_din <= x"005f0e89";
		wait for Clk_period;
		Addr <=  "00001110100010";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00001110100011";
		Trees_din <= x"ff690f3d";
		wait for Clk_period;
		Addr <=  "00001110100100";
		Trees_din <= x"0307f528";
		wait for Clk_period;
		Addr <=  "00001110100101";
		Trees_din <= x"18003308";
		wait for Clk_period;
		Addr <=  "00001110100110";
		Trees_din <= x"0b046404";
		wait for Clk_period;
		Addr <=  "00001110100111";
		Trees_din <= x"ff700f3d";
		wait for Clk_period;
		Addr <=  "00001110101000";
		Trees_din <= x"ffe90f3d";
		wait for Clk_period;
		Addr <=  "00001110101001";
		Trees_din <= x"1900a910";
		wait for Clk_period;
		Addr <=  "00001110101010";
		Trees_din <= x"07005508";
		wait for Clk_period;
		Addr <=  "00001110101011";
		Trees_din <= x"0b062504";
		wait for Clk_period;
		Addr <=  "00001110101100";
		Trees_din <= x"ff950f3d";
		wait for Clk_period;
		Addr <=  "00001110101101";
		Trees_din <= x"004f0f3d";
		wait for Clk_period;
		Addr <=  "00001110101110";
		Trees_din <= x"09005604";
		wait for Clk_period;
		Addr <=  "00001110101111";
		Trees_din <= x"00240f3d";
		wait for Clk_period;
		Addr <=  "00001110110000";
		Trees_din <= x"ffd20f3d";
		wait for Clk_period;
		Addr <=  "00001110110001";
		Trees_din <= x"17006c08";
		wait for Clk_period;
		Addr <=  "00001110110010";
		Trees_din <= x"14011b04";
		wait for Clk_period;
		Addr <=  "00001110110011";
		Trees_din <= x"002b0f3d";
		wait for Clk_period;
		Addr <=  "00001110110100";
		Trees_din <= x"ff910f3d";
		wait for Clk_period;
		Addr <=  "00001110110101";
		Trees_din <= x"0afcbf04";
		wait for Clk_period;
		Addr <=  "00001110110110";
		Trees_din <= x"00030f3d";
		wait for Clk_period;
		Addr <=  "00001110110111";
		Trees_din <= x"00ba0f3d";
		wait for Clk_period;
		Addr <=  "00001110111000";
		Trees_din <= x"0e03c01c";
		wait for Clk_period;
		Addr <=  "00001110111001";
		Trees_din <= x"05fde510";
		wait for Clk_period;
		Addr <=  "00001110111010";
		Trees_din <= x"12020c08";
		wait for Clk_period;
		Addr <=  "00001110111011";
		Trees_din <= x"0c015d04";
		wait for Clk_period;
		Addr <=  "00001110111100";
		Trees_din <= x"fff70f3d";
		wait for Clk_period;
		Addr <=  "00001110111101";
		Trees_din <= x"00520f3d";
		wait for Clk_period;
		Addr <=  "00001110111110";
		Trees_din <= x"00f8f604";
		wait for Clk_period;
		Addr <=  "00001110111111";
		Trees_din <= x"000c0f3d";
		wait for Clk_period;
		Addr <=  "00001111000000";
		Trees_din <= x"00960f3d";
		wait for Clk_period;
		Addr <=  "00001111000001";
		Trees_din <= x"0b028608";
		wait for Clk_period;
		Addr <=  "00001111000010";
		Trees_din <= x"11007904";
		wait for Clk_period;
		Addr <=  "00001111000011";
		Trees_din <= x"fff40f3d";
		wait for Clk_period;
		Addr <=  "00001111000100";
		Trees_din <= x"ff240f3d";
		wait for Clk_period;
		Addr <=  "00001111000101";
		Trees_din <= x"00920f3d";
		wait for Clk_period;
		Addr <=  "00001111000110";
		Trees_din <= x"0c020308";
		wait for Clk_period;
		Addr <=  "00001111000111";
		Trees_din <= x"030a7404";
		wait for Clk_period;
		Addr <=  "00001111001000";
		Trees_din <= x"ffa10f3d";
		wait for Clk_period;
		Addr <=  "00001111001001";
		Trees_din <= x"00800f3d";
		wait for Clk_period;
		Addr <=  "00001111001010";
		Trees_din <= x"06f53904";
		wait for Clk_period;
		Addr <=  "00001111001011";
		Trees_din <= x"ff410f3d";
		wait for Clk_period;
		Addr <=  "00001111001100";
		Trees_din <= x"04050404";
		wait for Clk_period;
		Addr <=  "00001111001101";
		Trees_din <= x"006c0f3d";
		wait for Clk_period;
		Addr <=  "00001111001110";
		Trees_din <= x"ff9c0f3d";
		wait for Clk_period;
		Addr <=  "00001111001111";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00001111010000";
		Trees_din <= x"ff690fe1";
		wait for Clk_period;
		Addr <=  "00001111010001";
		Trees_din <= x"0304d328";
		wait for Clk_period;
		Addr <=  "00001111010010";
		Trees_din <= x"0403b018";
		wait for Clk_period;
		Addr <=  "00001111010011";
		Trees_din <= x"06fa4510";
		wait for Clk_period;
		Addr <=  "00001111010100";
		Trees_din <= x"0f019c08";
		wait for Clk_period;
		Addr <=  "00001111010101";
		Trees_din <= x"06f78904";
		wait for Clk_period;
		Addr <=  "00001111010110";
		Trees_din <= x"000c0fe1";
		wait for Clk_period;
		Addr <=  "00001111010111";
		Trees_din <= x"00a10fe1";
		wait for Clk_period;
		Addr <=  "00001111011000";
		Trees_din <= x"010b7604";
		wait for Clk_period;
		Addr <=  "00001111011001";
		Trees_din <= x"ff9c0fe1";
		wait for Clk_period;
		Addr <=  "00001111011010";
		Trees_din <= x"007e0fe1";
		wait for Clk_period;
		Addr <=  "00001111011011";
		Trees_din <= x"0efd0504";
		wait for Clk_period;
		Addr <=  "00001111011100";
		Trees_din <= x"ffe90fe1";
		wait for Clk_period;
		Addr <=  "00001111011101";
		Trees_din <= x"ff7b0fe1";
		wait for Clk_period;
		Addr <=  "00001111011110";
		Trees_din <= x"0ef9a904";
		wait for Clk_period;
		Addr <=  "00001111011111";
		Trees_din <= x"005c0fe1";
		wait for Clk_period;
		Addr <=  "00001111100000";
		Trees_din <= x"10059708";
		wait for Clk_period;
		Addr <=  "00001111100001";
		Trees_din <= x"09004a04";
		wait for Clk_period;
		Addr <=  "00001111100010";
		Trees_din <= x"fffc0fe1";
		wait for Clk_period;
		Addr <=  "00001111100011";
		Trees_din <= x"ff680fe1";
		wait for Clk_period;
		Addr <=  "00001111100100";
		Trees_din <= x"00310fe1";
		wait for Clk_period;
		Addr <=  "00001111100101";
		Trees_din <= x"030fb41c";
		wait for Clk_period;
		Addr <=  "00001111100110";
		Trees_din <= x"09004c0c";
		wait for Clk_period;
		Addr <=  "00001111100111";
		Trees_din <= x"1500b208";
		wait for Clk_period;
		Addr <=  "00001111101000";
		Trees_din <= x"01fa4c04";
		wait for Clk_period;
		Addr <=  "00001111101001";
		Trees_din <= x"ffec0fe1";
		wait for Clk_period;
		Addr <=  "00001111101010";
		Trees_din <= x"00800fe1";
		wait for Clk_period;
		Addr <=  "00001111101011";
		Trees_din <= x"ffda0fe1";
		wait for Clk_period;
		Addr <=  "00001111101100";
		Trees_din <= x"06f5ff08";
		wait for Clk_period;
		Addr <=  "00001111101101";
		Trees_din <= x"03075d04";
		wait for Clk_period;
		Addr <=  "00001111101110";
		Trees_din <= x"ff850fe1";
		wait for Clk_period;
		Addr <=  "00001111101111";
		Trees_din <= x"fff60fe1";
		wait for Clk_period;
		Addr <=  "00001111110000";
		Trees_din <= x"1603d704";
		wait for Clk_period;
		Addr <=  "00001111110001";
		Trees_din <= x"003a0fe1";
		wait for Clk_period;
		Addr <=  "00001111110010";
		Trees_din <= x"ffc80fe1";
		wait for Clk_period;
		Addr <=  "00001111110011";
		Trees_din <= x"00f79208";
		wait for Clk_period;
		Addr <=  "00001111110100";
		Trees_din <= x"09005704";
		wait for Clk_period;
		Addr <=  "00001111110101";
		Trees_din <= x"005f0fe1";
		wait for Clk_period;
		Addr <=  "00001111110110";
		Trees_din <= x"ffa00fe1";
		wait for Clk_period;
		Addr <=  "00001111110111";
		Trees_din <= x"008d0fe1";
		wait for Clk_period;
		Addr <=  "00001111111000";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00001111111001";
		Trees_din <= x"ff6a1075";
		wait for Clk_period;
		Addr <=  "00001111111010";
		Trees_din <= x"030fb43c";
		wait for Clk_period;
		Addr <=  "00001111111011";
		Trees_din <= x"1100a220";
		wait for Clk_period;
		Addr <=  "00001111111100";
		Trees_din <= x"16021810";
		wait for Clk_period;
		Addr <=  "00001111111101";
		Trees_din <= x"09005408";
		wait for Clk_period;
		Addr <=  "00001111111110";
		Trees_din <= x"12fdea04";
		wait for Clk_period;
		Addr <=  "00001111111111";
		Trees_din <= x"ffcc1075";
		wait for Clk_period;
		Addr <=  "00010000000000";
		Trees_din <= x"006a1075";
		wait for Clk_period;
		Addr <=  "00010000000001";
		Trees_din <= x"03096504";
		wait for Clk_period;
		Addr <=  "00010000000010";
		Trees_din <= x"ff7d1075";
		wait for Clk_period;
		Addr <=  "00010000000011";
		Trees_din <= x"00131075";
		wait for Clk_period;
		Addr <=  "00010000000100";
		Trees_din <= x"06f54908";
		wait for Clk_period;
		Addr <=  "00010000000101";
		Trees_din <= x"07005704";
		wait for Clk_period;
		Addr <=  "00010000000110";
		Trees_din <= x"ff9c1075";
		wait for Clk_period;
		Addr <=  "00010000000111";
		Trees_din <= x"003e1075";
		wait for Clk_period;
		Addr <=  "00010000001000";
		Trees_din <= x"0a04b804";
		wait for Clk_period;
		Addr <=  "00010000001001";
		Trees_din <= x"006e1075";
		wait for Clk_period;
		Addr <=  "00010000001010";
		Trees_din <= x"ffab1075";
		wait for Clk_period;
		Addr <=  "00010000001011";
		Trees_din <= x"0303820c";
		wait for Clk_period;
		Addr <=  "00010000001100";
		Trees_din <= x"1603fe08";
		wait for Clk_period;
		Addr <=  "00010000001101";
		Trees_din <= x"08000904";
		wait for Clk_period;
		Addr <=  "00010000001110";
		Trees_din <= x"002d1075";
		wait for Clk_period;
		Addr <=  "00010000001111";
		Trees_din <= x"ff891075";
		wait for Clk_period;
		Addr <=  "00010000010000";
		Trees_din <= x"00701075";
		wait for Clk_period;
		Addr <=  "00010000010001";
		Trees_din <= x"01feb608";
		wait for Clk_period;
		Addr <=  "00010000010010";
		Trees_din <= x"01fbee04";
		wait for Clk_period;
		Addr <=  "00010000010011";
		Trees_din <= x"00141075";
		wait for Clk_period;
		Addr <=  "00010000010100";
		Trees_din <= x"ffc51075";
		wait for Clk_period;
		Addr <=  "00010000010101";
		Trees_din <= x"16011204";
		wait for Clk_period;
		Addr <=  "00010000010110";
		Trees_din <= x"006c1075";
		wait for Clk_period;
		Addr <=  "00010000010111";
		Trees_din <= x"00081075";
		wait for Clk_period;
		Addr <=  "00010000011000";
		Trees_din <= x"08002508";
		wait for Clk_period;
		Addr <=  "00010000011001";
		Trees_din <= x"09005704";
		wait for Clk_period;
		Addr <=  "00010000011010";
		Trees_din <= x"00591075";
		wait for Clk_period;
		Addr <=  "00010000011011";
		Trees_din <= x"ffa61075";
		wait for Clk_period;
		Addr <=  "00010000011100";
		Trees_din <= x"008a1075";
		wait for Clk_period;
		Addr <=  "00010000011101";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00010000011110";
		Trees_din <= x"ff6b10f1";
		wait for Clk_period;
		Addr <=  "00010000011111";
		Trees_din <= x"0308a91c";
		wait for Clk_period;
		Addr <=  "00010000100000";
		Trees_din <= x"05f86604";
		wait for Clk_period;
		Addr <=  "00010000100001";
		Trees_din <= x"ff7d10f1";
		wait for Clk_period;
		Addr <=  "00010000100010";
		Trees_din <= x"18003308";
		wait for Clk_period;
		Addr <=  "00010000100011";
		Trees_din <= x"0b043104";
		wait for Clk_period;
		Addr <=  "00010000100100";
		Trees_din <= x"ff7610f1";
		wait for Clk_period;
		Addr <=  "00010000100101";
		Trees_din <= x"000710f1";
		wait for Clk_period;
		Addr <=  "00010000100110";
		Trees_din <= x"09005808";
		wait for Clk_period;
		Addr <=  "00010000100111";
		Trees_din <= x"0101df04";
		wait for Clk_period;
		Addr <=  "00010000101000";
		Trees_din <= x"ffef10f1";
		wait for Clk_period;
		Addr <=  "00010000101001";
		Trees_din <= x"003f10f1";
		wait for Clk_period;
		Addr <=  "00010000101010";
		Trees_din <= x"0e023004";
		wait for Clk_period;
		Addr <=  "00010000101011";
		Trees_din <= x"ff9c10f1";
		wait for Clk_period;
		Addr <=  "00010000101100";
		Trees_din <= x"001b10f1";
		wait for Clk_period;
		Addr <=  "00010000101101";
		Trees_din <= x"18003708";
		wait for Clk_period;
		Addr <=  "00010000101110";
		Trees_din <= x"0a029104";
		wait for Clk_period;
		Addr <=  "00010000101111";
		Trees_din <= x"009310f1";
		wait for Clk_period;
		Addr <=  "00010000110000";
		Trees_din <= x"001a10f1";
		wait for Clk_period;
		Addr <=  "00010000110001";
		Trees_din <= x"18003808";
		wait for Clk_period;
		Addr <=  "00010000110010";
		Trees_din <= x"0d023404";
		wait for Clk_period;
		Addr <=  "00010000110011";
		Trees_din <= x"001f10f1";
		wait for Clk_period;
		Addr <=  "00010000110100";
		Trees_din <= x"ff3f10f1";
		wait for Clk_period;
		Addr <=  "00010000110101";
		Trees_din <= x"04041b08";
		wait for Clk_period;
		Addr <=  "00010000110110";
		Trees_din <= x"1603f104";
		wait for Clk_period;
		Addr <=  "00010000110111";
		Trees_din <= x"007410f1";
		wait for Clk_period;
		Addr <=  "00010000111000";
		Trees_din <= x"fff210f1";
		wait for Clk_period;
		Addr <=  "00010000111001";
		Trees_din <= x"02001704";
		wait for Clk_period;
		Addr <=  "00010000111010";
		Trees_din <= x"002310f1";
		wait for Clk_period;
		Addr <=  "00010000111011";
		Trees_din <= x"ffb710f1";
		wait for Clk_period;
		Addr <=  "00010000111100";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00010000111101";
		Trees_din <= x"ff6c1155";
		wait for Clk_period;
		Addr <=  "00010000111110";
		Trees_din <= x"030fb424";
		wait for Clk_period;
		Addr <=  "00010000111111";
		Trees_din <= x"02091320";
		wait for Clk_period;
		Addr <=  "00010001000000";
		Trees_din <= x"1100a210";
		wait for Clk_period;
		Addr <=  "00010001000001";
		Trees_din <= x"1a00c908";
		wait for Clk_period;
		Addr <=  "00010001000010";
		Trees_din <= x"14018a04";
		wait for Clk_period;
		Addr <=  "00010001000011";
		Trees_din <= x"002d1155";
		wait for Clk_period;
		Addr <=  "00010001000100";
		Trees_din <= x"ffa81155";
		wait for Clk_period;
		Addr <=  "00010001000101";
		Trees_din <= x"0802ea04";
		wait for Clk_period;
		Addr <=  "00010001000110";
		Trees_din <= x"00681155";
		wait for Clk_period;
		Addr <=  "00010001000111";
		Trees_din <= x"ffc51155";
		wait for Clk_period;
		Addr <=  "00010001001000";
		Trees_din <= x"03038208";
		wait for Clk_period;
		Addr <=  "00010001001001";
		Trees_din <= x"05fac804";
		wait for Clk_period;
		Addr <=  "00010001001010";
		Trees_din <= x"00111155";
		wait for Clk_period;
		Addr <=  "00010001001011";
		Trees_din <= x"ff921155";
		wait for Clk_period;
		Addr <=  "00010001001100";
		Trees_din <= x"01feb604";
		wait for Clk_period;
		Addr <=  "00010001001101";
		Trees_din <= x"ffe71155";
		wait for Clk_period;
		Addr <=  "00010001001110";
		Trees_din <= x"00271155";
		wait for Clk_period;
		Addr <=  "00010001001111";
		Trees_din <= x"ff8e1155";
		wait for Clk_period;
		Addr <=  "00010001010000";
		Trees_din <= x"10055008";
		wait for Clk_period;
		Addr <=  "00010001010001";
		Trees_din <= x"1b004804";
		wait for Clk_period;
		Addr <=  "00010001010010";
		Trees_din <= x"00831155";
		wait for Clk_period;
		Addr <=  "00010001010011";
		Trees_din <= x"00201155";
		wait for Clk_period;
		Addr <=  "00010001010100";
		Trees_din <= x"ffdf1155";
		wait for Clk_period;
		Addr <=  "00010001010101";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00010001010110";
		Trees_din <= x"ff6e1211";
		wait for Clk_period;
		Addr <=  "00010001010111";
		Trees_din <= x"030bbf34";
		wait for Clk_period;
		Addr <=  "00010001011000";
		Trees_din <= x"1f000120";
		wait for Clk_period;
		Addr <=  "00010001011001";
		Trees_din <= x"00050810";
		wait for Clk_period;
		Addr <=  "00010001011010";
		Trees_din <= x"00019008";
		wait for Clk_period;
		Addr <=  "00010001011011";
		Trees_din <= x"0c01d804";
		wait for Clk_period;
		Addr <=  "00010001011100";
		Trees_din <= x"00131211";
		wait for Clk_period;
		Addr <=  "00010001011101";
		Trees_din <= x"ffd01211";
		wait for Clk_period;
		Addr <=  "00010001011110";
		Trees_din <= x"02fe5a04";
		wait for Clk_period;
		Addr <=  "00010001011111";
		Trees_din <= x"00151211";
		wait for Clk_period;
		Addr <=  "00010001100000";
		Trees_din <= x"ff821211";
		wait for Clk_period;
		Addr <=  "00010001100001";
		Trees_din <= x"0007fa08";
		wait for Clk_period;
		Addr <=  "00010001100010";
		Trees_din <= x"15009b04";
		wait for Clk_period;
		Addr <=  "00010001100011";
		Trees_din <= x"ffd31211";
		wait for Clk_period;
		Addr <=  "00010001100100";
		Trees_din <= x"00af1211";
		wait for Clk_period;
		Addr <=  "00010001100101";
		Trees_din <= x"0e03d504";
		wait for Clk_period;
		Addr <=  "00010001100110";
		Trees_din <= x"ff8c1211";
		wait for Clk_period;
		Addr <=  "00010001100111";
		Trees_din <= x"00671211";
		wait for Clk_period;
		Addr <=  "00010001101000";
		Trees_din <= x"0700550c";
		wait for Clk_period;
		Addr <=  "00010001101001";
		Trees_din <= x"10faf604";
		wait for Clk_period;
		Addr <=  "00010001101010";
		Trees_din <= x"00601211";
		wait for Clk_period;
		Addr <=  "00010001101011";
		Trees_din <= x"1a010704";
		wait for Clk_period;
		Addr <=  "00010001101100";
		Trees_din <= x"ff831211";
		wait for Clk_period;
		Addr <=  "00010001101101";
		Trees_din <= x"00151211";
		wait for Clk_period;
		Addr <=  "00010001101110";
		Trees_din <= x"0002d304";
		wait for Clk_period;
		Addr <=  "00010001101111";
		Trees_din <= x"00971211";
		wait for Clk_period;
		Addr <=  "00010001110000";
		Trees_din <= x"00161211";
		wait for Clk_period;
		Addr <=  "00010001110001";
		Trees_din <= x"19009b14";
		wait for Clk_period;
		Addr <=  "00010001110010";
		Trees_din <= x"0bfb7a0c";
		wait for Clk_period;
		Addr <=  "00010001110011";
		Trees_din <= x"0f028e08";
		wait for Clk_period;
		Addr <=  "00010001110100";
		Trees_din <= x"13ff8c04";
		wait for Clk_period;
		Addr <=  "00010001110101";
		Trees_din <= x"fff01211";
		wait for Clk_period;
		Addr <=  "00010001110110";
		Trees_din <= x"006d1211";
		wait for Clk_period;
		Addr <=  "00010001110111";
		Trees_din <= x"ffab1211";
		wait for Clk_period;
		Addr <=  "00010001111000";
		Trees_din <= x"1b004704";
		wait for Clk_period;
		Addr <=  "00010001111001";
		Trees_din <= x"00881211";
		wait for Clk_period;
		Addr <=  "00010001111010";
		Trees_din <= x"00111211";
		wait for Clk_period;
		Addr <=  "00010001111011";
		Trees_din <= x"0f012b10";
		wait for Clk_period;
		Addr <=  "00010001111100";
		Trees_din <= x"1e005d08";
		wait for Clk_period;
		Addr <=  "00010001111101";
		Trees_din <= x"13ffb104";
		wait for Clk_period;
		Addr <=  "00010001111110";
		Trees_din <= x"006f1211";
		wait for Clk_period;
		Addr <=  "00010001111111";
		Trees_din <= x"ffd11211";
		wait for Clk_period;
		Addr <=  "00010010000000";
		Trees_din <= x"1400b104";
		wait for Clk_period;
		Addr <=  "00010010000001";
		Trees_din <= x"ffd21211";
		wait for Clk_period;
		Addr <=  "00010010000010";
		Trees_din <= x"ff6c1211";
		wait for Clk_period;
		Addr <=  "00010010000011";
		Trees_din <= x"00671211";
		wait for Clk_period;
		Addr <=  "00010010000100";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00010010000101";
		Trees_din <= x"ff6f12ed";
		wait for Clk_period;
		Addr <=  "00010010000110";
		Trees_din <= x"0305c734";
		wait for Clk_period;
		Addr <=  "00010010000111";
		Trees_din <= x"00060120";
		wait for Clk_period;
		Addr <=  "00010010001000";
		Trees_din <= x"0c01bf10";
		wait for Clk_period;
		Addr <=  "00010010001001";
		Trees_din <= x"1b004708";
		wait for Clk_period;
		Addr <=  "00010010001010";
		Trees_din <= x"12fe8304";
		wait for Clk_period;
		Addr <=  "00010010001011";
		Trees_din <= x"003412ed";
		wait for Clk_period;
		Addr <=  "00010010001100";
		Trees_din <= x"ffc012ed";
		wait for Clk_period;
		Addr <=  "00010010001101";
		Trees_din <= x"11018f04";
		wait for Clk_period;
		Addr <=  "00010010001110";
		Trees_din <= x"ffff12ed";
		wait for Clk_period;
		Addr <=  "00010010001111";
		Trees_din <= x"007912ed";
		wait for Clk_period;
		Addr <=  "00010010010000";
		Trees_din <= x"20040008";
		wait for Clk_period;
		Addr <=  "00010010010001";
		Trees_din <= x"17000404";
		wait for Clk_period;
		Addr <=  "00010010010010";
		Trees_din <= x"ffe512ed";
		wait for Clk_period;
		Addr <=  "00010010010011";
		Trees_din <= x"005112ed";
		wait for Clk_period;
		Addr <=  "00010010010100";
		Trees_din <= x"07005b04";
		wait for Clk_period;
		Addr <=  "00010010010101";
		Trees_din <= x"ff6912ed";
		wait for Clk_period;
		Addr <=  "00010010010110";
		Trees_din <= x"ffed12ed";
		wait for Clk_period;
		Addr <=  "00010010010111";
		Trees_din <= x"0007fa08";
		wait for Clk_period;
		Addr <=  "00010010011000";
		Trees_din <= x"15009b04";
		wait for Clk_period;
		Addr <=  "00010010011001";
		Trees_din <= x"ffe912ed";
		wait for Clk_period;
		Addr <=  "00010010011010";
		Trees_din <= x"00db12ed";
		wait for Clk_period;
		Addr <=  "00010010011011";
		Trees_din <= x"03038208";
		wait for Clk_period;
		Addr <=  "00010010011100";
		Trees_din <= x"14007804";
		wait for Clk_period;
		Addr <=  "00010010011101";
		Trees_din <= x"fffe12ed";
		wait for Clk_period;
		Addr <=  "00010010011110";
		Trees_din <= x"ff8312ed";
		wait for Clk_period;
		Addr <=  "00010010011111";
		Trees_din <= x"003b12ed";
		wait for Clk_period;
		Addr <=  "00010010100000";
		Trees_din <= x"0c015d18";
		wait for Clk_period;
		Addr <=  "00010010100001";
		Trees_din <= x"07005008";
		wait for Clk_period;
		Addr <=  "00010010100010";
		Trees_din <= x"06f52304";
		wait for Clk_period;
		Addr <=  "00010010100011";
		Trees_din <= x"002312ed";
		wait for Clk_period;
		Addr <=  "00010010100100";
		Trees_din <= x"008212ed";
		wait for Clk_period;
		Addr <=  "00010010100101";
		Trees_din <= x"030b0208";
		wait for Clk_period;
		Addr <=  "00010010100110";
		Trees_din <= x"02fb4704";
		wait for Clk_period;
		Addr <=  "00010010100111";
		Trees_din <= x"006212ed";
		wait for Clk_period;
		Addr <=  "00010010101000";
		Trees_din <= x"ffb112ed";
		wait for Clk_period;
		Addr <=  "00010010101001";
		Trees_din <= x"12020704";
		wait for Clk_period;
		Addr <=  "00010010101010";
		Trees_din <= x"fff912ed";
		wait for Clk_period;
		Addr <=  "00010010101011";
		Trees_din <= x"008112ed";
		wait for Clk_period;
		Addr <=  "00010010101100";
		Trees_din <= x"06f3df10";
		wait for Clk_period;
		Addr <=  "00010010101101";
		Trees_din <= x"0c02fd08";
		wait for Clk_period;
		Addr <=  "00010010101110";
		Trees_din <= x"02000604";
		wait for Clk_period;
		Addr <=  "00010010101111";
		Trees_din <= x"ffee12ed";
		wait for Clk_period;
		Addr <=  "00010010110000";
		Trees_din <= x"ff7512ed";
		wait for Clk_period;
		Addr <=  "00010010110001";
		Trees_din <= x"09005604";
		wait for Clk_period;
		Addr <=  "00010010110010";
		Trees_din <= x"005b12ed";
		wait for Clk_period;
		Addr <=  "00010010110011";
		Trees_din <= x"ffc912ed";
		wait for Clk_period;
		Addr <=  "00010010110100";
		Trees_din <= x"02fbdf08";
		wait for Clk_period;
		Addr <=  "00010010110101";
		Trees_din <= x"1a00bf04";
		wait for Clk_period;
		Addr <=  "00010010110110";
		Trees_din <= x"004d12ed";
		wait for Clk_period;
		Addr <=  "00010010110111";
		Trees_din <= x"ffb012ed";
		wait for Clk_period;
		Addr <=  "00010010111000";
		Trees_din <= x"09005204";
		wait for Clk_period;
		Addr <=  "00010010111001";
		Trees_din <= x"001112ed";
		wait for Clk_period;
		Addr <=  "00010010111010";
		Trees_din <= x"006f12ed";
		wait for Clk_period;
		Addr <=  "00010010111011";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00010010111100";
		Trees_din <= x"ff711341";
		wait for Clk_period;
		Addr <=  "00010010111101";
		Trees_din <= x"04f85504";
		wait for Clk_period;
		Addr <=  "00010010111110";
		Trees_din <= x"ff9b1341";
		wait for Clk_period;
		Addr <=  "00010010111111";
		Trees_din <= x"02091320";
		wait for Clk_period;
		Addr <=  "00010011000000";
		Trees_din <= x"04041b10";
		wait for Clk_period;
		Addr <=  "00010011000001";
		Trees_din <= x"09005308";
		wait for Clk_period;
		Addr <=  "00010011000010";
		Trees_din <= x"0afc7c04";
		wait for Clk_period;
		Addr <=  "00010011000011";
		Trees_din <= x"ffbb1341";
		wait for Clk_period;
		Addr <=  "00010011000100";
		Trees_din <= x"00281341";
		wait for Clk_period;
		Addr <=  "00010011000101";
		Trees_din <= x"06f96104";
		wait for Clk_period;
		Addr <=  "00010011000110";
		Trees_din <= x"005b1341";
		wait for Clk_period;
		Addr <=  "00010011000111";
		Trees_din <= x"ffee1341";
		wait for Clk_period;
		Addr <=  "00010011001000";
		Trees_din <= x"0304d308";
		wait for Clk_period;
		Addr <=  "00010011001001";
		Trees_din <= x"0ef9a904";
		wait for Clk_period;
		Addr <=  "00010011001010";
		Trees_din <= x"00581341";
		wait for Clk_period;
		Addr <=  "00010011001011";
		Trees_din <= x"ffa01341";
		wait for Clk_period;
		Addr <=  "00010011001100";
		Trees_din <= x"09004f04";
		wait for Clk_period;
		Addr <=  "00010011001101";
		Trees_din <= x"00621341";
		wait for Clk_period;
		Addr <=  "00010011001110";
		Trees_din <= x"fff81341";
		wait for Clk_period;
		Addr <=  "00010011001111";
		Trees_din <= x"ff981341";
		wait for Clk_period;
		Addr <=  "00010011010000";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00010011010001";
		Trees_din <= x"ff72142d";
		wait for Clk_period;
		Addr <=  "00010011010010";
		Trees_din <= x"0308a93c";
		wait for Clk_period;
		Addr <=  "00010011010011";
		Trees_din <= x"0800c71c";
		wait for Clk_period;
		Addr <=  "00010011010100";
		Trees_din <= x"08009110";
		wait for Clk_period;
		Addr <=  "00010011010101";
		Trees_din <= x"0101fc08";
		wait for Clk_period;
		Addr <=  "00010011010110";
		Trees_din <= x"09005704";
		wait for Clk_period;
		Addr <=  "00010011010111";
		Trees_din <= x"ff92142d";
		wait for Clk_period;
		Addr <=  "00010011011000";
		Trees_din <= x"001a142d";
		wait for Clk_period;
		Addr <=  "00010011011001";
		Trees_din <= x"0200f004";
		wait for Clk_period;
		Addr <=  "00010011011010";
		Trees_din <= x"ffde142d";
		wait for Clk_period;
		Addr <=  "00010011011011";
		Trees_din <= x"005d142d";
		wait for Clk_period;
		Addr <=  "00010011011100";
		Trees_din <= x"0302da04";
		wait for Clk_period;
		Addr <=  "00010011011101";
		Trees_din <= x"ffa6142d";
		wait for Clk_period;
		Addr <=  "00010011011110";
		Trees_din <= x"04fe5b04";
		wait for Clk_period;
		Addr <=  "00010011011111";
		Trees_din <= x"000b142d";
		wait for Clk_period;
		Addr <=  "00010011100000";
		Trees_din <= x"00a4142d";
		wait for Clk_period;
		Addr <=  "00010011100001";
		Trees_din <= x"0801f410";
		wait for Clk_period;
		Addr <=  "00010011100010";
		Trees_din <= x"0d004408";
		wait for Clk_period;
		Addr <=  "00010011100011";
		Trees_din <= x"10fbe004";
		wait for Clk_period;
		Addr <=  "00010011100100";
		Trees_din <= x"0054142d";
		wait for Clk_period;
		Addr <=  "00010011100101";
		Trees_din <= x"ffd4142d";
		wait for Clk_period;
		Addr <=  "00010011100110";
		Trees_din <= x"0307f504";
		wait for Clk_period;
		Addr <=  "00010011100111";
		Trees_din <= x"ff73142d";
		wait for Clk_period;
		Addr <=  "00010011101000";
		Trees_din <= x"fff4142d";
		wait for Clk_period;
		Addr <=  "00010011101001";
		Trees_din <= x"07005808";
		wait for Clk_period;
		Addr <=  "00010011101010";
		Trees_din <= x"17016004";
		wait for Clk_period;
		Addr <=  "00010011101011";
		Trees_din <= x"ffb4142d";
		wait for Clk_period;
		Addr <=  "00010011101100";
		Trees_din <= x"003d142d";
		wait for Clk_period;
		Addr <=  "00010011101101";
		Trees_din <= x"11028604";
		wait for Clk_period;
		Addr <=  "00010011101110";
		Trees_din <= x"fffa142d";
		wait for Clk_period;
		Addr <=  "00010011101111";
		Trees_din <= x"009f142d";
		wait for Clk_period;
		Addr <=  "00010011110000";
		Trees_din <= x"01fdeb20";
		wait for Clk_period;
		Addr <=  "00010011110001";
		Trees_din <= x"01fd0910";
		wait for Clk_period;
		Addr <=  "00010011110010";
		Trees_din <= x"05fde508";
		wait for Clk_period;
		Addr <=  "00010011110011";
		Trees_din <= x"09005404";
		wait for Clk_period;
		Addr <=  "00010011110100";
		Trees_din <= x"0063142d";
		wait for Clk_period;
		Addr <=  "00010011110101";
		Trees_din <= x"ffff142d";
		wait for Clk_period;
		Addr <=  "00010011110110";
		Trees_din <= x"0b028404";
		wait for Clk_period;
		Addr <=  "00010011110111";
		Trees_din <= x"ff60142d";
		wait for Clk_period;
		Addr <=  "00010011111000";
		Trees_din <= x"0060142d";
		wait for Clk_period;
		Addr <=  "00010011111001";
		Trees_din <= x"04041b08";
		wait for Clk_period;
		Addr <=  "00010011111010";
		Trees_din <= x"01fd4e04";
		wait for Clk_period;
		Addr <=  "00010011111011";
		Trees_din <= x"ffd0142d";
		wait for Clk_period;
		Addr <=  "00010011111100";
		Trees_din <= x"0042142d";
		wait for Clk_period;
		Addr <=  "00010011111101";
		Trees_din <= x"030bbf04";
		wait for Clk_period;
		Addr <=  "00010011111110";
		Trees_din <= x"ff65142d";
		wait for Clk_period;
		Addr <=  "00010011111111";
		Trees_din <= x"ffec142d";
		wait for Clk_period;
		Addr <=  "00010100000000";
		Trees_din <= x"0d02910c";
		wait for Clk_period;
		Addr <=  "00010100000001";
		Trees_din <= x"06f05e04";
		wait for Clk_period;
		Addr <=  "00010100000010";
		Trees_din <= x"0000142d";
		wait for Clk_period;
		Addr <=  "00010100000011";
		Trees_din <= x"08003e04";
		wait for Clk_period;
		Addr <=  "00010100000100";
		Trees_din <= x"001f142d";
		wait for Clk_period;
		Addr <=  "00010100000101";
		Trees_din <= x"008f142d";
		wait for Clk_period;
		Addr <=  "00010100000110";
		Trees_din <= x"16032808";
		wait for Clk_period;
		Addr <=  "00010100000111";
		Trees_din <= x"1d004604";
		wait for Clk_period;
		Addr <=  "00010100001000";
		Trees_din <= x"006f142d";
		wait for Clk_period;
		Addr <=  "00010100001001";
		Trees_din <= x"fff4142d";
		wait for Clk_period;
		Addr <=  "00010100001010";
		Trees_din <= x"ff9c142d";
		wait for Clk_period;
		Addr <=  "00010100001011";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00010100001100";
		Trees_din <= x"ff7514a1";
		wait for Clk_period;
		Addr <=  "00010100001101";
		Trees_din <= x"0008bf2c";
		wait for Clk_period;
		Addr <=  "00010100001110";
		Trees_din <= x"0006341c";
		wait for Clk_period;
		Addr <=  "00010100001111";
		Trees_din <= x"0301f90c";
		wait for Clk_period;
		Addr <=  "00010100010000";
		Trees_din <= x"1d004b04";
		wait for Clk_period;
		Addr <=  "00010100010001";
		Trees_din <= x"ff7f14a1";
		wait for Clk_period;
		Addr <=  "00010100010010";
		Trees_din <= x"0e025204";
		wait for Clk_period;
		Addr <=  "00010100010011";
		Trees_din <= x"ffdb14a1";
		wait for Clk_period;
		Addr <=  "00010100010100";
		Trees_din <= x"005414a1";
		wait for Clk_period;
		Addr <=  "00010100010101";
		Trees_din <= x"09004c08";
		wait for Clk_period;
		Addr <=  "00010100010110";
		Trees_din <= x"1500b204";
		wait for Clk_period;
		Addr <=  "00010100010111";
		Trees_din <= x"005714a1";
		wait for Clk_period;
		Addr <=  "00010100011000";
		Trees_din <= x"ffe214a1";
		wait for Clk_period;
		Addr <=  "00010100011001";
		Trees_din <= x"01020f04";
		wait for Clk_period;
		Addr <=  "00010100011010";
		Trees_din <= x"ffef14a1";
		wait for Clk_period;
		Addr <=  "00010100011011";
		Trees_din <= x"002314a1";
		wait for Clk_period;
		Addr <=  "00010100011100";
		Trees_din <= x"1800420c";
		wait for Clk_period;
		Addr <=  "00010100011101";
		Trees_din <= x"0c02bd08";
		wait for Clk_period;
		Addr <=  "00010100011110";
		Trees_din <= x"06f61f04";
		wait for Clk_period;
		Addr <=  "00010100011111";
		Trees_din <= x"003414a1";
		wait for Clk_period;
		Addr <=  "00010100100000";
		Trees_din <= x"00bf14a1";
		wait for Clk_period;
		Addr <=  "00010100100001";
		Trees_din <= x"000814a1";
		wait for Clk_period;
		Addr <=  "00010100100010";
		Trees_din <= x"ffd014a1";
		wait for Clk_period;
		Addr <=  "00010100100011";
		Trees_din <= x"18004204";
		wait for Clk_period;
		Addr <=  "00010100100100";
		Trees_din <= x"ff8414a1";
		wait for Clk_period;
		Addr <=  "00010100100101";
		Trees_din <= x"1a00bd04";
		wait for Clk_period;
		Addr <=  "00010100100110";
		Trees_din <= x"ffad14a1";
		wait for Clk_period;
		Addr <=  "00010100100111";
		Trees_din <= x"007c14a1";
		wait for Clk_period;
		Addr <=  "00010100101000";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00010100101001";
		Trees_din <= x"ff771565";
		wait for Clk_period;
		Addr <=  "00010100101010";
		Trees_din <= x"030bbf34";
		wait for Clk_period;
		Addr <=  "00010100101011";
		Trees_din <= x"06f5231c";
		wait for Clk_period;
		Addr <=  "00010100101100";
		Trees_din <= x"0f00a310";
		wait for Clk_period;
		Addr <=  "00010100101101";
		Trees_din <= x"0b040e08";
		wait for Clk_period;
		Addr <=  "00010100101110";
		Trees_din <= x"1a00fc04";
		wait for Clk_period;
		Addr <=  "00010100101111";
		Trees_din <= x"00541565";
		wait for Clk_period;
		Addr <=  "00010100110000";
		Trees_din <= x"ffc61565";
		wait for Clk_period;
		Addr <=  "00010100110001";
		Trees_din <= x"18004204";
		wait for Clk_period;
		Addr <=  "00010100110010";
		Trees_din <= x"ff841565";
		wait for Clk_period;
		Addr <=  "00010100110011";
		Trees_din <= x"001d1565";
		wait for Clk_period;
		Addr <=  "00010100110100";
		Trees_din <= x"1203b708";
		wait for Clk_period;
		Addr <=  "00010100110101";
		Trees_din <= x"13f92e04";
		wait for Clk_period;
		Addr <=  "00010100110110";
		Trees_din <= x"00211565";
		wait for Clk_period;
		Addr <=  "00010100110111";
		Trees_din <= x"ff7b1565";
		wait for Clk_period;
		Addr <=  "00010100111000";
		Trees_din <= x"00391565";
		wait for Clk_period;
		Addr <=  "00010100111001";
		Trees_din <= x"06f56508";
		wait for Clk_period;
		Addr <=  "00010100111010";
		Trees_din <= x"18004404";
		wait for Clk_period;
		Addr <=  "00010100111011";
		Trees_din <= x"00b61565";
		wait for Clk_period;
		Addr <=  "00010100111100";
		Trees_din <= x"ffd71565";
		wait for Clk_period;
		Addr <=  "00010100111101";
		Trees_din <= x"07005b08";
		wait for Clk_period;
		Addr <=  "00010100111110";
		Trees_din <= x"0b045004";
		wait for Clk_period;
		Addr <=  "00010100111111";
		Trees_din <= x"ffda1565";
		wait for Clk_period;
		Addr <=  "00010101000000";
		Trees_din <= x"00201565";
		wait for Clk_period;
		Addr <=  "00010101000001";
		Trees_din <= x"0d030504";
		wait for Clk_period;
		Addr <=  "00010101000010";
		Trees_din <= x"00671565";
		wait for Clk_period;
		Addr <=  "00010101000011";
		Trees_din <= x"ffda1565";
		wait for Clk_period;
		Addr <=  "00010101000100";
		Trees_din <= x"1500a51c";
		wait for Clk_period;
		Addr <=  "00010101000101";
		Trees_din <= x"0408ca0c";
		wait for Clk_period;
		Addr <=  "00010101000110";
		Trees_din <= x"14003908";
		wait for Clk_period;
		Addr <=  "00010101000111";
		Trees_din <= x"13fdca04";
		wait for Clk_period;
		Addr <=  "00010101001000";
		Trees_din <= x"00431565";
		wait for Clk_period;
		Addr <=  "00010101001001";
		Trees_din <= x"ffc01565";
		wait for Clk_period;
		Addr <=  "00010101001010";
		Trees_din <= x"00891565";
		wait for Clk_period;
		Addr <=  "00010101001011";
		Trees_din <= x"11028408";
		wait for Clk_period;
		Addr <=  "00010101001100";
		Trees_din <= x"08007804";
		wait for Clk_period;
		Addr <=  "00010101001101";
		Trees_din <= x"ffd91565";
		wait for Clk_period;
		Addr <=  "00010101001110";
		Trees_din <= x"00601565";
		wait for Clk_period;
		Addr <=  "00010101001111";
		Trees_din <= x"13ff8c04";
		wait for Clk_period;
		Addr <=  "00010101010000";
		Trees_din <= x"ffa11565";
		wait for Clk_period;
		Addr <=  "00010101010001";
		Trees_din <= x"00081565";
		wait for Clk_period;
		Addr <=  "00010101010010";
		Trees_din <= x"1701c508";
		wait for Clk_period;
		Addr <=  "00010101010011";
		Trees_din <= x"11028304";
		wait for Clk_period;
		Addr <=  "00010101010100";
		Trees_din <= x"00601565";
		wait for Clk_period;
		Addr <=  "00010101010101";
		Trees_din <= x"ffe21565";
		wait for Clk_period;
		Addr <=  "00010101010110";
		Trees_din <= x"0b04c704";
		wait for Clk_period;
		Addr <=  "00010101010111";
		Trees_din <= x"fffa1565";
		wait for Clk_period;
		Addr <=  "00010101011000";
		Trees_din <= x"ff851565";
		wait for Clk_period;
		Addr <=  "00010101011001";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00010101011010";
		Trees_din <= x"ff791629";
		wait for Clk_period;
		Addr <=  "00010101011011";
		Trees_din <= x"03075d28";
		wait for Clk_period;
		Addr <=  "00010101011100";
		Trees_din <= x"10fa2808";
		wait for Clk_period;
		Addr <=  "00010101011101";
		Trees_din <= x"08000b04";
		wait for Clk_period;
		Addr <=  "00010101011110";
		Trees_din <= x"001d1629";
		wait for Clk_period;
		Addr <=  "00010101011111";
		Trees_din <= x"ff7b1629";
		wait for Clk_period;
		Addr <=  "00010101100000";
		Trees_din <= x"09005610";
		wait for Clk_period;
		Addr <=  "00010101100001";
		Trees_din <= x"1500a908";
		wait for Clk_period;
		Addr <=  "00010101100010";
		Trees_din <= x"11fea004";
		wait for Clk_period;
		Addr <=  "00010101100011";
		Trees_din <= x"ffb11629";
		wait for Clk_period;
		Addr <=  "00010101100100";
		Trees_din <= x"003c1629";
		wait for Clk_period;
		Addr <=  "00010101100101";
		Trees_din <= x"06fad804";
		wait for Clk_period;
		Addr <=  "00010101100110";
		Trees_din <= x"ff8f1629";
		wait for Clk_period;
		Addr <=  "00010101100111";
		Trees_din <= x"00271629";
		wait for Clk_period;
		Addr <=  "00010101101000";
		Trees_din <= x"08021408";
		wait for Clk_period;
		Addr <=  "00010101101001";
		Trees_din <= x"08002104";
		wait for Clk_period;
		Addr <=  "00010101101010";
		Trees_din <= x"00091629";
		wait for Clk_period;
		Addr <=  "00010101101011";
		Trees_din <= x"ff721629";
		wait for Clk_period;
		Addr <=  "00010101101100";
		Trees_din <= x"0f00f204";
		wait for Clk_period;
		Addr <=  "00010101101101";
		Trees_din <= x"00681629";
		wait for Clk_period;
		Addr <=  "00010101101110";
		Trees_din <= x"ff9d1629";
		wait for Clk_period;
		Addr <=  "00010101101111";
		Trees_din <= x"0bfb1c1c";
		wait for Clk_period;
		Addr <=  "00010101110000";
		Trees_din <= x"05fbb610";
		wait for Clk_period;
		Addr <=  "00010101110001";
		Trees_din <= x"03096508";
		wait for Clk_period;
		Addr <=  "00010101110010";
		Trees_din <= x"0afb1504";
		wait for Clk_period;
		Addr <=  "00010101110011";
		Trees_din <= x"00171629";
		wait for Clk_period;
		Addr <=  "00010101110100";
		Trees_din <= x"ff961629";
		wait for Clk_period;
		Addr <=  "00010101110101";
		Trees_din <= x"02018704";
		wait for Clk_period;
		Addr <=  "00010101110110";
		Trees_din <= x"007d1629";
		wait for Clk_period;
		Addr <=  "00010101110111";
		Trees_din <= x"ffd51629";
		wait for Clk_period;
		Addr <=  "00010101111000";
		Trees_din <= x"0d025404";
		wait for Clk_period;
		Addr <=  "00010101111001";
		Trees_din <= x"ff731629";
		wait for Clk_period;
		Addr <=  "00010101111010";
		Trees_din <= x"1b003304";
		wait for Clk_period;
		Addr <=  "00010101111011";
		Trees_din <= x"ffb91629";
		wait for Clk_period;
		Addr <=  "00010101111100";
		Trees_din <= x"00431629";
		wait for Clk_period;
		Addr <=  "00010101111101";
		Trees_din <= x"06f3b40c";
		wait for Clk_period;
		Addr <=  "00010101111110";
		Trees_din <= x"11027d08";
		wait for Clk_period;
		Addr <=  "00010101111111";
		Trees_din <= x"1c003304";
		wait for Clk_period;
		Addr <=  "00010110000000";
		Trees_din <= x"ffc41629";
		wait for Clk_period;
		Addr <=  "00010110000001";
		Trees_din <= x"00551629";
		wait for Clk_period;
		Addr <=  "00010110000010";
		Trees_din <= x"ff8a1629";
		wait for Clk_period;
		Addr <=  "00010110000011";
		Trees_din <= x"0afadb08";
		wait for Clk_period;
		Addr <=  "00010110000100";
		Trees_din <= x"0c008104";
		wait for Clk_period;
		Addr <=  "00010110000101";
		Trees_din <= x"ffb91629";
		wait for Clk_period;
		Addr <=  "00010110000110";
		Trees_din <= x"00351629";
		wait for Clk_period;
		Addr <=  "00010110000111";
		Trees_din <= x"01fa9904";
		wait for Clk_period;
		Addr <=  "00010110001000";
		Trees_din <= x"fffa1629";
		wait for Clk_period;
		Addr <=  "00010110001001";
		Trees_din <= x"006a1629";
		wait for Clk_period;
		Addr <=  "00010110001010";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00010110001011";
		Trees_din <= x"ff7c16ed";
		wait for Clk_period;
		Addr <=  "00010110001100";
		Trees_din <= x"0308a924";
		wait for Clk_period;
		Addr <=  "00010110001101";
		Trees_din <= x"05f86604";
		wait for Clk_period;
		Addr <=  "00010110001110";
		Trees_din <= x"ff8c16ed";
		wait for Clk_period;
		Addr <=  "00010110001111";
		Trees_din <= x"0800c710";
		wait for Clk_period;
		Addr <=  "00010110010000";
		Trees_din <= x"08009108";
		wait for Clk_period;
		Addr <=  "00010110010001";
		Trees_din <= x"0101fc04";
		wait for Clk_period;
		Addr <=  "00010110010010";
		Trees_din <= x"ffcb16ed";
		wait for Clk_period;
		Addr <=  "00010110010011";
		Trees_din <= x"002c16ed";
		wait for Clk_period;
		Addr <=  "00010110010100";
		Trees_din <= x"04014904";
		wait for Clk_period;
		Addr <=  "00010110010101";
		Trees_din <= x"000816ed";
		wait for Clk_period;
		Addr <=  "00010110010110";
		Trees_din <= x"008416ed";
		wait for Clk_period;
		Addr <=  "00010110010111";
		Trees_din <= x"0801f408";
		wait for Clk_period;
		Addr <=  "00010110011000";
		Trees_din <= x"03075d04";
		wait for Clk_period;
		Addr <=  "00010110011001";
		Trees_din <= x"ff8a16ed";
		wait for Clk_period;
		Addr <=  "00010110011010";
		Trees_din <= x"000616ed";
		wait for Clk_period;
		Addr <=  "00010110011011";
		Trees_din <= x"11028804";
		wait for Clk_period;
		Addr <=  "00010110011100";
		Trees_din <= x"ffeb16ed";
		wait for Clk_period;
		Addr <=  "00010110011101";
		Trees_din <= x"005d16ed";
		wait for Clk_period;
		Addr <=  "00010110011110";
		Trees_din <= x"1b003b20";
		wait for Clk_period;
		Addr <=  "00010110011111";
		Trees_din <= x"1900a610";
		wait for Clk_period;
		Addr <=  "00010110100000";
		Trees_din <= x"0e03c008";
		wait for Clk_period;
		Addr <=  "00010110100001";
		Trees_din <= x"00011804";
		wait for Clk_period;
		Addr <=  "00010110100010";
		Trees_din <= x"007e16ed";
		wait for Clk_period;
		Addr <=  "00010110100011";
		Trees_din <= x"001116ed";
		wait for Clk_period;
		Addr <=  "00010110100100";
		Trees_din <= x"02fc9504";
		wait for Clk_period;
		Addr <=  "00010110100101";
		Trees_din <= x"ffb516ed";
		wait for Clk_period;
		Addr <=  "00010110100110";
		Trees_din <= x"002916ed";
		wait for Clk_period;
		Addr <=  "00010110100111";
		Trees_din <= x"1d003b08";
		wait for Clk_period;
		Addr <=  "00010110101000";
		Trees_din <= x"0b04cb04";
		wait for Clk_period;
		Addr <=  "00010110101001";
		Trees_din <= x"005616ed";
		wait for Clk_period;
		Addr <=  "00010110101010";
		Trees_din <= x"ffd916ed";
		wait for Clk_period;
		Addr <=  "00010110101011";
		Trees_din <= x"16033104";
		wait for Clk_period;
		Addr <=  "00010110101100";
		Trees_din <= x"fff316ed";
		wait for Clk_period;
		Addr <=  "00010110101101";
		Trees_din <= x"ff6716ed";
		wait for Clk_period;
		Addr <=  "00010110101110";
		Trees_din <= x"19008a0c";
		wait for Clk_period;
		Addr <=  "00010110101111";
		Trees_din <= x"1403d008";
		wait for Clk_period;
		Addr <=  "00010110110000";
		Trees_din <= x"08002504";
		wait for Clk_period;
		Addr <=  "00010110110001";
		Trees_din <= x"fff316ed";
		wait for Clk_period;
		Addr <=  "00010110110010";
		Trees_din <= x"007216ed";
		wait for Clk_period;
		Addr <=  "00010110110011";
		Trees_din <= x"ffc116ed";
		wait for Clk_period;
		Addr <=  "00010110110100";
		Trees_din <= x"07005908";
		wait for Clk_period;
		Addr <=  "00010110110101";
		Trees_din <= x"030bbf04";
		wait for Clk_period;
		Addr <=  "00010110110110";
		Trees_din <= x"ff8016ed";
		wait for Clk_period;
		Addr <=  "00010110110111";
		Trees_din <= x"000416ed";
		wait for Clk_period;
		Addr <=  "00010110111000";
		Trees_din <= x"09005704";
		wait for Clk_period;
		Addr <=  "00010110111001";
		Trees_din <= x"ffd816ed";
		wait for Clk_period;
		Addr <=  "00010110111010";
		Trees_din <= x"005916ed";
		wait for Clk_period;
		Addr <=  "00010110111011";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00010110111100";
		Trees_din <= x"ff7e1779";
		wait for Clk_period;
		Addr <=  "00010110111101";
		Trees_din <= x"20040020";
		wait for Clk_period;
		Addr <=  "00010110111110";
		Trees_din <= x"0f03fc1c";
		wait for Clk_period;
		Addr <=  "00010110111111";
		Trees_din <= x"11028310";
		wait for Clk_period;
		Addr <=  "00010111000000";
		Trees_din <= x"13fa6408";
		wait for Clk_period;
		Addr <=  "00010111000001";
		Trees_din <= x"0d017e04";
		wait for Clk_period;
		Addr <=  "00010111000010";
		Trees_din <= x"003b1779";
		wait for Clk_period;
		Addr <=  "00010111000011";
		Trees_din <= x"ffb61779";
		wait for Clk_period;
		Addr <=  "00010111000100";
		Trees_din <= x"07005a04";
		wait for Clk_period;
		Addr <=  "00010111000101";
		Trees_din <= x"00881779";
		wait for Clk_period;
		Addr <=  "00010111000110";
		Trees_din <= x"00091779";
		wait for Clk_period;
		Addr <=  "00010111000111";
		Trees_din <= x"18004204";
		wait for Clk_period;
		Addr <=  "00010111001000";
		Trees_din <= x"ffa51779";
		wait for Clk_period;
		Addr <=  "00010111001001";
		Trees_din <= x"0306c204";
		wait for Clk_period;
		Addr <=  "00010111001010";
		Trees_din <= x"ffdb1779";
		wait for Clk_period;
		Addr <=  "00010111001011";
		Trees_din <= x"006c1779";
		wait for Clk_period;
		Addr <=  "00010111001100";
		Trees_din <= x"ffb31779";
		wait for Clk_period;
		Addr <=  "00010111001101";
		Trees_din <= x"01f8ef04";
		wait for Clk_period;
		Addr <=  "00010111001110";
		Trees_din <= x"00641779";
		wait for Clk_period;
		Addr <=  "00010111001111";
		Trees_din <= x"1c003810";
		wait for Clk_period;
		Addr <=  "00010111010000";
		Trees_din <= x"1c003508";
		wait for Clk_period;
		Addr <=  "00010111010001";
		Trees_din <= x"1102cd04";
		wait for Clk_period;
		Addr <=  "00010111010010";
		Trees_din <= x"ffe91779";
		wait for Clk_period;
		Addr <=  "00010111010011";
		Trees_din <= x"002b1779";
		wait for Clk_period;
		Addr <=  "00010111010100";
		Trees_din <= x"17000104";
		wait for Clk_period;
		Addr <=  "00010111010101";
		Trees_din <= x"ffea1779";
		wait for Clk_period;
		Addr <=  "00010111010110";
		Trees_din <= x"00851779";
		wait for Clk_period;
		Addr <=  "00010111010111";
		Trees_din <= x"01030e08";
		wait for Clk_period;
		Addr <=  "00010111011000";
		Trees_din <= x"02ff0f04";
		wait for Clk_period;
		Addr <=  "00010111011001";
		Trees_din <= x"fff81779";
		wait for Clk_period;
		Addr <=  "00010111011010";
		Trees_din <= x"ffa21779";
		wait for Clk_period;
		Addr <=  "00010111011011";
		Trees_din <= x"01070104";
		wait for Clk_period;
		Addr <=  "00010111011100";
		Trees_din <= x"00411779";
		wait for Clk_period;
		Addr <=  "00010111011101";
		Trees_din <= x"ffc71779";
		wait for Clk_period;
		Addr <=  "00010111011110";
		Trees_din <= x"000b1e34";
		wait for Clk_period;
		Addr <=  "00010111011111";
		Trees_din <= x"02091330";
		wait for Clk_period;
		Addr <=  "00010111100000";
		Trees_din <= x"04041b14";
		wait for Clk_period;
		Addr <=  "00010111100001";
		Trees_din <= x"04f85504";
		wait for Clk_period;
		Addr <=  "00010111100010";
		Trees_din <= x"ffaf17e5";
		wait for Clk_period;
		Addr <=  "00010111100011";
		Trees_din <= x"0bf94d08";
		wait for Clk_period;
		Addr <=  "00010111100100";
		Trees_din <= x"1004ad04";
		wait for Clk_period;
		Addr <=  "00010111100101";
		Trees_din <= x"002917e5";
		wait for Clk_period;
		Addr <=  "00010111100110";
		Trees_din <= x"ff9717e5";
		wait for Clk_period;
		Addr <=  "00010111100111";
		Trees_din <= x"16006d04";
		wait for Clk_period;
		Addr <=  "00010111101000";
		Trees_din <= x"ffe417e5";
		wait for Clk_period;
		Addr <=  "00010111101001";
		Trees_din <= x"002d17e5";
		wait for Clk_period;
		Addr <=  "00010111101010";
		Trees_din <= x"02fece0c";
		wait for Clk_period;
		Addr <=  "00010111101011";
		Trees_din <= x"0e03d008";
		wait for Clk_period;
		Addr <=  "00010111101100";
		Trees_din <= x"1c003804";
		wait for Clk_period;
		Addr <=  "00010111101101";
		Trees_din <= x"003f17e5";
		wait for Clk_period;
		Addr <=  "00010111101110";
		Trees_din <= x"ffed17e5";
		wait for Clk_period;
		Addr <=  "00010111101111";
		Trees_din <= x"ffb017e5";
		wait for Clk_period;
		Addr <=  "00010111110000";
		Trees_din <= x"00feee08";
		wait for Clk_period;
		Addr <=  "00010111110001";
		Trees_din <= x"09005704";
		wait for Clk_period;
		Addr <=  "00010111110010";
		Trees_din <= x"001817e5";
		wait for Clk_period;
		Addr <=  "00010111110011";
		Trees_din <= x"ffb717e5";
		wait for Clk_period;
		Addr <=  "00010111110100";
		Trees_din <= x"0c026d04";
		wait for Clk_period;
		Addr <=  "00010111110101";
		Trees_din <= x"ff7517e5";
		wait for Clk_period;
		Addr <=  "00010111110110";
		Trees_din <= x"000217e5";
		wait for Clk_period;
		Addr <=  "00010111110111";
		Trees_din <= x"ff9817e5";
		wait for Clk_period;
		Addr <=  "00010111111000";
		Trees_din <= x"ff8117e5";
		wait for Clk_period;
		Addr <=  "00010111111001";
		Trees_din <= x"0302911c";
		wait for Clk_period;
		Addr <=  "00010111111010";
		Trees_din <= x"1b002d08";
		wait for Clk_period;
		Addr <=  "00010111111011";
		Trees_din <= x"18003804";
		wait for Clk_period;
		Addr <=  "00010111111100";
		Trees_din <= x"ffac18a9";
		wait for Clk_period;
		Addr <=  "00010111111101";
		Trees_din <= x"008b18a9";
		wait for Clk_period;
		Addr <=  "00010111111110";
		Trees_din <= x"07005e10";
		wait for Clk_period;
		Addr <=  "00010111111111";
		Trees_din <= x"2100000c";
		wait for Clk_period;
		Addr <=  "00011000000000";
		Trees_din <= x"08000908";
		wait for Clk_period;
		Addr <=  "00011000000001";
		Trees_din <= x"12023a04";
		wait for Clk_period;
		Addr <=  "00011000000010";
		Trees_din <= x"ffae18a9";
		wait for Clk_period;
		Addr <=  "00011000000011";
		Trees_din <= x"003218a9";
		wait for Clk_period;
		Addr <=  "00011000000100";
		Trees_din <= x"ff7c18a9";
		wait for Clk_period;
		Addr <=  "00011000000101";
		Trees_din <= x"001d18a9";
		wait for Clk_period;
		Addr <=  "00011000000110";
		Trees_din <= x"001c18a9";
		wait for Clk_period;
		Addr <=  "00011000000111";
		Trees_din <= x"09004c14";
		wait for Clk_period;
		Addr <=  "00011000001000";
		Trees_din <= x"0002570c";
		wait for Clk_period;
		Addr <=  "00011000001001";
		Trees_din <= x"01021f08";
		wait for Clk_period;
		Addr <=  "00011000001010";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00011000001011";
		Trees_din <= x"000b18a9";
		wait for Clk_period;
		Addr <=  "00011000001100";
		Trees_din <= x"007e18a9";
		wait for Clk_period;
		Addr <=  "00011000001101";
		Trees_din <= x"fffe18a9";
		wait for Clk_period;
		Addr <=  "00011000001110";
		Trees_din <= x"0c006e04";
		wait for Clk_period;
		Addr <=  "00011000001111";
		Trees_din <= x"005d18a9";
		wait for Clk_period;
		Addr <=  "00011000010000";
		Trees_din <= x"ffac18a9";
		wait for Clk_period;
		Addr <=  "00011000010001";
		Trees_din <= x"09005114";
		wait for Clk_period;
		Addr <=  "00011000010010";
		Trees_din <= x"07005108";
		wait for Clk_period;
		Addr <=  "00011000010011";
		Trees_din <= x"0c021604";
		wait for Clk_period;
		Addr <=  "00011000010100";
		Trees_din <= x"007118a9";
		wait for Clk_period;
		Addr <=  "00011000010101";
		Trees_din <= x"ffba18a9";
		wait for Clk_period;
		Addr <=  "00011000010110";
		Trees_din <= x"06f48704";
		wait for Clk_period;
		Addr <=  "00011000010111";
		Trees_din <= x"000e18a9";
		wait for Clk_period;
		Addr <=  "00011000011000";
		Trees_din <= x"0d030d04";
		wait for Clk_period;
		Addr <=  "00011000011001";
		Trees_din <= x"ff7b18a9";
		wait for Clk_period;
		Addr <=  "00011000011010";
		Trees_din <= x"ffe218a9";
		wait for Clk_period;
		Addr <=  "00011000011011";
		Trees_din <= x"1400c110";
		wait for Clk_period;
		Addr <=  "00011000011100";
		Trees_din <= x"0afae408";
		wait for Clk_period;
		Addr <=  "00011000011101";
		Trees_din <= x"0af78704";
		wait for Clk_period;
		Addr <=  "00011000011110";
		Trees_din <= x"000218a9";
		wait for Clk_period;
		Addr <=  "00011000011111";
		Trees_din <= x"ff9a18a9";
		wait for Clk_period;
		Addr <=  "00011000100000";
		Trees_din <= x"0308a904";
		wait for Clk_period;
		Addr <=  "00011000100001";
		Trees_din <= x"ffdf18a9";
		wait for Clk_period;
		Addr <=  "00011000100010";
		Trees_din <= x"003718a9";
		wait for Clk_period;
		Addr <=  "00011000100011";
		Trees_din <= x"0afca708";
		wait for Clk_period;
		Addr <=  "00011000100100";
		Trees_din <= x"02034a04";
		wait for Clk_period;
		Addr <=  "00011000100101";
		Trees_din <= x"005718a9";
		wait for Clk_period;
		Addr <=  "00011000100110";
		Trees_din <= x"ffdb18a9";
		wait for Clk_period;
		Addr <=  "00011000100111";
		Trees_din <= x"02ff0b04";
		wait for Clk_period;
		Addr <=  "00011000101000";
		Trees_din <= x"001e18a9";
		wait for Clk_period;
		Addr <=  "00011000101001";
		Trees_din <= x"ffdc18a9";
		wait for Clk_period;
		Addr <=  "00011000101010";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00011000101011";
		Trees_din <= x"ff87195d";
		wait for Clk_period;
		Addr <=  "00011000101100";
		Trees_din <= x"030a7430";
		wait for Clk_period;
		Addr <=  "00011000101101";
		Trees_din <= x"00fba514";
		wait for Clk_period;
		Addr <=  "00011000101110";
		Trees_din <= x"1d003a08";
		wait for Clk_period;
		Addr <=  "00011000101111";
		Trees_din <= x"1b002b04";
		wait for Clk_period;
		Addr <=  "00011000110000";
		Trees_din <= x"ffb6195d";
		wait for Clk_period;
		Addr <=  "00011000110001";
		Trees_din <= x"0065195d";
		wait for Clk_period;
		Addr <=  "00011000110010";
		Trees_din <= x"08000004";
		wait for Clk_period;
		Addr <=  "00011000110011";
		Trees_din <= x"0024195d";
		wait for Clk_period;
		Addr <=  "00011000110100";
		Trees_din <= x"04004504";
		wait for Clk_period;
		Addr <=  "00011000110101";
		Trees_din <= x"fff6195d";
		wait for Clk_period;
		Addr <=  "00011000110110";
		Trees_din <= x"ff89195d";
		wait for Clk_period;
		Addr <=  "00011000110111";
		Trees_din <= x"16006d0c";
		wait for Clk_period;
		Addr <=  "00011000111000";
		Trees_din <= x"02ffb908";
		wait for Clk_period;
		Addr <=  "00011000111001";
		Trees_din <= x"1b003404";
		wait for Clk_period;
		Addr <=  "00011000111010";
		Trees_din <= x"005d195d";
		wait for Clk_period;
		Addr <=  "00011000111011";
		Trees_din <= x"ffde195d";
		wait for Clk_period;
		Addr <=  "00011000111100";
		Trees_din <= x"ff7f195d";
		wait for Clk_period;
		Addr <=  "00011000111101";
		Trees_din <= x"09005408";
		wait for Clk_period;
		Addr <=  "00011000111110";
		Trees_din <= x"05ff4a04";
		wait for Clk_period;
		Addr <=  "00011000111111";
		Trees_din <= x"ffdd195d";
		wait for Clk_period;
		Addr <=  "00011001000000";
		Trees_din <= x"0055195d";
		wait for Clk_period;
		Addr <=  "00011001000001";
		Trees_din <= x"06f42b04";
		wait for Clk_period;
		Addr <=  "00011001000010";
		Trees_din <= x"ffc8195d";
		wait for Clk_period;
		Addr <=  "00011001000011";
		Trees_din <= x"003f195d";
		wait for Clk_period;
		Addr <=  "00011001000100";
		Trees_din <= x"0d01f714";
		wait for Clk_period;
		Addr <=  "00011001000101";
		Trees_din <= x"1a00a108";
		wait for Clk_period;
		Addr <=  "00011001000110";
		Trees_din <= x"0f006104";
		wait for Clk_period;
		Addr <=  "00011001000111";
		Trees_din <= x"0016195d";
		wait for Clk_period;
		Addr <=  "00011001001000";
		Trees_din <= x"ffba195d";
		wait for Clk_period;
		Addr <=  "00011001001001";
		Trees_din <= x"02fd1508";
		wait for Clk_period;
		Addr <=  "00011001001010";
		Trees_din <= x"0f007b04";
		wait for Clk_period;
		Addr <=  "00011001001011";
		Trees_din <= x"ffe6195d";
		wait for Clk_period;
		Addr <=  "00011001001100";
		Trees_din <= x"004a195d";
		wait for Clk_period;
		Addr <=  "00011001001101";
		Trees_din <= x"007f195d";
		wait for Clk_period;
		Addr <=  "00011001001110";
		Trees_din <= x"15009008";
		wait for Clk_period;
		Addr <=  "00011001001111";
		Trees_din <= x"0f003f04";
		wait for Clk_period;
		Addr <=  "00011001010000";
		Trees_din <= x"ffee195d";
		wait for Clk_period;
		Addr <=  "00011001010001";
		Trees_din <= x"0071195d";
		wait for Clk_period;
		Addr <=  "00011001010010";
		Trees_din <= x"13012a08";
		wait for Clk_period;
		Addr <=  "00011001010011";
		Trees_din <= x"1d003b04";
		wait for Clk_period;
		Addr <=  "00011001010100";
		Trees_din <= x"0014195d";
		wait for Clk_period;
		Addr <=  "00011001010101";
		Trees_din <= x"ffa6195d";
		wait for Clk_period;
		Addr <=  "00011001010110";
		Trees_din <= x"0057195d";
		wait for Clk_period;
		Addr <=  "00011001010111";
		Trees_din <= x"000b1e64";
		wait for Clk_period;
		Addr <=  "00011001011000";
		Trees_din <= x"0308a93c";
		wait for Clk_period;
		Addr <=  "00011001011001";
		Trees_din <= x"0800c71c";
		wait for Clk_period;
		Addr <=  "00011001011010";
		Trees_din <= x"08009110";
		wait for Clk_period;
		Addr <=  "00011001011011";
		Trees_din <= x"0400ad08";
		wait for Clk_period;
		Addr <=  "00011001011100";
		Trees_din <= x"04fdef04";
		wait for Clk_period;
		Addr <=  "00011001011101";
		Trees_din <= x"ffd61a29";
		wait for Clk_period;
		Addr <=  "00011001011110";
		Trees_din <= x"00601a29";
		wait for Clk_period;
		Addr <=  "00011001011111";
		Trees_din <= x"08000104";
		wait for Clk_period;
		Addr <=  "00011001100000";
		Trees_din <= x"00361a29";
		wait for Clk_period;
		Addr <=  "00011001100001";
		Trees_din <= x"ffc21a29";
		wait for Clk_period;
		Addr <=  "00011001100010";
		Trees_din <= x"06f55004";
		wait for Clk_period;
		Addr <=  "00011001100011";
		Trees_din <= x"fffc1a29";
		wait for Clk_period;
		Addr <=  "00011001100100";
		Trees_din <= x"04022404";
		wait for Clk_period;
		Addr <=  "00011001100101";
		Trees_din <= x"00101a29";
		wait for Clk_period;
		Addr <=  "00011001100110";
		Trees_din <= x"008b1a29";
		wait for Clk_period;
		Addr <=  "00011001100111";
		Trees_din <= x"0801f410";
		wait for Clk_period;
		Addr <=  "00011001101000";
		Trees_din <= x"0d004408";
		wait for Clk_period;
		Addr <=  "00011001101001";
		Trees_din <= x"0e002904";
		wait for Clk_period;
		Addr <=  "00011001101010";
		Trees_din <= x"ffe21a29";
		wait for Clk_period;
		Addr <=  "00011001101011";
		Trees_din <= x"003b1a29";
		wait for Clk_period;
		Addr <=  "00011001101100";
		Trees_din <= x"0307f504";
		wait for Clk_period;
		Addr <=  "00011001101101";
		Trees_din <= x"ff831a29";
		wait for Clk_period;
		Addr <=  "00011001101110";
		Trees_din <= x"fffa1a29";
		wait for Clk_period;
		Addr <=  "00011001101111";
		Trees_din <= x"07005808";
		wait for Clk_period;
		Addr <=  "00011001110000";
		Trees_din <= x"11009a04";
		wait for Clk_period;
		Addr <=  "00011001110001";
		Trees_din <= x"00211a29";
		wait for Clk_period;
		Addr <=  "00011001110010";
		Trees_din <= x"ffb01a29";
		wait for Clk_period;
		Addr <=  "00011001110011";
		Trees_din <= x"0b028704";
		wait for Clk_period;
		Addr <=  "00011001110100";
		Trees_din <= x"006a1a29";
		wait for Clk_period;
		Addr <=  "00011001110101";
		Trees_din <= x"ffd81a29";
		wait for Clk_period;
		Addr <=  "00011001110110";
		Trees_din <= x"01fdeb18";
		wait for Clk_period;
		Addr <=  "00011001110111";
		Trees_din <= x"01fd0910";
		wait for Clk_period;
		Addr <=  "00011001111000";
		Trees_din <= x"1004f608";
		wait for Clk_period;
		Addr <=  "00011001111001";
		Trees_din <= x"1a00d204";
		wait for Clk_period;
		Addr <=  "00011001111010";
		Trees_din <= x"00071a29";
		wait for Clk_period;
		Addr <=  "00011001111011";
		Trees_din <= x"006b1a29";
		wait for Clk_period;
		Addr <=  "00011001111100";
		Trees_din <= x"0c014004";
		wait for Clk_period;
		Addr <=  "00011001111101";
		Trees_din <= x"ffa31a29";
		wait for Clk_period;
		Addr <=  "00011001111110";
		Trees_din <= x"00341a29";
		wait for Clk_period;
		Addr <=  "00011001111111";
		Trees_din <= x"04041b04";
		wait for Clk_period;
		Addr <=  "00011010000000";
		Trees_din <= x"00101a29";
		wait for Clk_period;
		Addr <=  "00011010000001";
		Trees_din <= x"ff9f1a29";
		wait for Clk_period;
		Addr <=  "00011010000010";
		Trees_din <= x"07005204";
		wait for Clk_period;
		Addr <=  "00011010000011";
		Trees_din <= x"ffe61a29";
		wait for Clk_period;
		Addr <=  "00011010000100";
		Trees_din <= x"0afaf204";
		wait for Clk_period;
		Addr <=  "00011010000101";
		Trees_din <= x"00011a29";
		wait for Clk_period;
		Addr <=  "00011010000110";
		Trees_din <= x"06f3ec04";
		wait for Clk_period;
		Addr <=  "00011010000111";
		Trees_din <= x"00241a29";
		wait for Clk_period;
		Addr <=  "00011010001000";
		Trees_din <= x"00831a29";
		wait for Clk_period;
		Addr <=  "00011010001001";
		Trees_din <= x"ff891a29";
		wait for Clk_period;
		Addr <=  "00011010001010";
		Trees_din <= x"000b1e40";
		wait for Clk_period;
		Addr <=  "00011010001011";
		Trees_din <= x"1500b138";
		wait for Clk_period;
		Addr <=  "00011010001100";
		Trees_din <= x"030bbf1c";
		wait for Clk_period;
		Addr <=  "00011010001101";
		Trees_din <= x"1f000110";
		wait for Clk_period;
		Addr <=  "00011010001110";
		Trees_din <= x"00050808";
		wait for Clk_period;
		Addr <=  "00011010001111";
		Trees_din <= x"00019004";
		wait for Clk_period;
		Addr <=  "00011010010000";
		Trees_din <= x"fffb1aad";
		wait for Clk_period;
		Addr <=  "00011010010001";
		Trees_din <= x"ffb81aad";
		wait for Clk_period;
		Addr <=  "00011010010010";
		Trees_din <= x"15009704";
		wait for Clk_period;
		Addr <=  "00011010010011";
		Trees_din <= x"ffc91aad";
		wait for Clk_period;
		Addr <=  "00011010010100";
		Trees_din <= x"00581aad";
		wait for Clk_period;
		Addr <=  "00011010010101";
		Trees_din <= x"22000004";
		wait for Clk_period;
		Addr <=  "00011010010110";
		Trees_din <= x"00621aad";
		wait for Clk_period;
		Addr <=  "00011010010111";
		Trees_din <= x"0a01e504";
		wait for Clk_period;
		Addr <=  "00011010011000";
		Trees_din <= x"ffc61aad";
		wait for Clk_period;
		Addr <=  "00011010011001";
		Trees_din <= x"00321aad";
		wait for Clk_period;
		Addr <=  "00011010011010";
		Trees_din <= x"09005710";
		wait for Clk_period;
		Addr <=  "00011010011011";
		Trees_din <= x"05fbbb08";
		wait for Clk_period;
		Addr <=  "00011010011100";
		Trees_din <= x"0409d604";
		wait for Clk_period;
		Addr <=  "00011010011101";
		Trees_din <= x"00721aad";
		wait for Clk_period;
		Addr <=  "00011010011110";
		Trees_din <= x"00171aad";
		wait for Clk_period;
		Addr <=  "00011010011111";
		Trees_din <= x"0bfb1c04";
		wait for Clk_period;
		Addr <=  "00011010100000";
		Trees_din <= x"ffc21aad";
		wait for Clk_period;
		Addr <=  "00011010100001";
		Trees_din <= x"00561aad";
		wait for Clk_period;
		Addr <=  "00011010100010";
		Trees_din <= x"09005704";
		wait for Clk_period;
		Addr <=  "00011010100011";
		Trees_din <= x"ffb01aad";
		wait for Clk_period;
		Addr <=  "00011010100100";
		Trees_din <= x"0f007b04";
		wait for Clk_period;
		Addr <=  "00011010100101";
		Trees_din <= x"fff61aad";
		wait for Clk_period;
		Addr <=  "00011010100110";
		Trees_din <= x"00531aad";
		wait for Clk_period;
		Addr <=  "00011010100111";
		Trees_din <= x"02fdc004";
		wait for Clk_period;
		Addr <=  "00011010101000";
		Trees_din <= x"00061aad";
		wait for Clk_period;
		Addr <=  "00011010101001";
		Trees_din <= x"ff971aad";
		wait for Clk_period;
		Addr <=  "00011010101010";
		Trees_din <= x"ff8d1aad";
		wait for Clk_period;
		Addr <=  "00011010101011";
		Trees_din <= x"0302911c";
		wait for Clk_period;
		Addr <=  "00011010101100";
		Trees_din <= x"06f7890c";
		wait for Clk_period;
		Addr <=  "00011010101101";
		Trees_din <= x"07005e08";
		wait for Clk_period;
		Addr <=  "00011010101110";
		Trees_din <= x"13014104";
		wait for Clk_period;
		Addr <=  "00011010101111";
		Trees_din <= x"ff7e1b81";
		wait for Clk_period;
		Addr <=  "00011010110000";
		Trees_din <= x"ffed1b81";
		wait for Clk_period;
		Addr <=  "00011010110001";
		Trees_din <= x"00241b81";
		wait for Clk_period;
		Addr <=  "00011010110010";
		Trees_din <= x"1700b204";
		wait for Clk_period;
		Addr <=  "00011010110011";
		Trees_din <= x"ff9d1b81";
		wait for Clk_period;
		Addr <=  "00011010110100";
		Trees_din <= x"0006ac08";
		wait for Clk_period;
		Addr <=  "00011010110101";
		Trees_din <= x"0005c704";
		wait for Clk_period;
		Addr <=  "00011010110110";
		Trees_din <= x"fff91b81";
		wait for Clk_period;
		Addr <=  "00011010110111";
		Trees_din <= x"008b1b81";
		wait for Clk_period;
		Addr <=  "00011010111000";
		Trees_din <= x"ffdf1b81";
		wait for Clk_period;
		Addr <=  "00011010111001";
		Trees_din <= x"0700592c";
		wait for Clk_period;
		Addr <=  "00011010111010";
		Trees_din <= x"17039720";
		wait for Clk_period;
		Addr <=  "00011010111011";
		Trees_din <= x"1b003a10";
		wait for Clk_period;
		Addr <=  "00011010111100";
		Trees_din <= x"18004208";
		wait for Clk_period;
		Addr <=  "00011010111101";
		Trees_din <= x"11017104";
		wait for Clk_period;
		Addr <=  "00011010111110";
		Trees_din <= x"001c1b81";
		wait for Clk_period;
		Addr <=  "00011010111111";
		Trees_din <= x"ffde1b81";
		wait for Clk_period;
		Addr <=  "00011011000000";
		Trees_din <= x"18004404";
		wait for Clk_period;
		Addr <=  "00011011000001";
		Trees_din <= x"00871b81";
		wait for Clk_period;
		Addr <=  "00011011000010";
		Trees_din <= x"ffed1b81";
		wait for Clk_period;
		Addr <=  "00011011000011";
		Trees_din <= x"19008408";
		wait for Clk_period;
		Addr <=  "00011011000100";
		Trees_din <= x"11018904";
		wait for Clk_period;
		Addr <=  "00011011000101";
		Trees_din <= x"ffcd1b81";
		wait for Clk_period;
		Addr <=  "00011011000110";
		Trees_din <= x"004e1b81";
		wait for Clk_period;
		Addr <=  "00011011000111";
		Trees_din <= x"030bbf04";
		wait for Clk_period;
		Addr <=  "00011011001000";
		Trees_din <= x"ff891b81";
		wait for Clk_period;
		Addr <=  "00011011001001";
		Trees_din <= x"00171b81";
		wait for Clk_period;
		Addr <=  "00011011001010";
		Trees_din <= x"05fb5604";
		wait for Clk_period;
		Addr <=  "00011011001011";
		Trees_din <= x"00701b81";
		wait for Clk_period;
		Addr <=  "00011011001100";
		Trees_din <= x"00fcaf04";
		wait for Clk_period;
		Addr <=  "00011011001101";
		Trees_din <= x"ffbd1b81";
		wait for Clk_period;
		Addr <=  "00011011001110";
		Trees_din <= x"00381b81";
		wait for Clk_period;
		Addr <=  "00011011001111";
		Trees_din <= x"00fa240c";
		wait for Clk_period;
		Addr <=  "00011011010000";
		Trees_din <= x"0f00a304";
		wait for Clk_period;
		Addr <=  "00011011010001";
		Trees_din <= x"002e1b81";
		wait for Clk_period;
		Addr <=  "00011011010010";
		Trees_din <= x"02ff0b04";
		wait for Clk_period;
		Addr <=  "00011011010011";
		Trees_din <= x"fff81b81";
		wait for Clk_period;
		Addr <=  "00011011010100";
		Trees_din <= x"ff9e1b81";
		wait for Clk_period;
		Addr <=  "00011011010101";
		Trees_din <= x"0306c20c";
		wait for Clk_period;
		Addr <=  "00011011010110";
		Trees_din <= x"19009808";
		wait for Clk_period;
		Addr <=  "00011011010111";
		Trees_din <= x"1c003b04";
		wait for Clk_period;
		Addr <=  "00011011011000";
		Trees_din <= x"00541b81";
		wait for Clk_period;
		Addr <=  "00011011011001";
		Trees_din <= x"fff01b81";
		wait for Clk_period;
		Addr <=  "00011011011010";
		Trees_din <= x"ff951b81";
		wait for Clk_period;
		Addr <=  "00011011011011";
		Trees_din <= x"14008008";
		wait for Clk_period;
		Addr <=  "00011011011100";
		Trees_din <= x"1100fa04";
		wait for Clk_period;
		Addr <=  "00011011011101";
		Trees_din <= x"00361b81";
		wait for Clk_period;
		Addr <=  "00011011011110";
		Trees_din <= x"ffd91b81";
		wait for Clk_period;
		Addr <=  "00011011011111";
		Trees_din <= x"007f1b81";
		wait for Clk_period;
		Addr <=  "00011011100000";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00011011100001";
		Trees_din <= x"0008bf44";
		wait for Clk_period;
		Addr <=  "00011011100010";
		Trees_din <= x"00063438";
		wait for Clk_period;
		Addr <=  "00011011100011";
		Trees_din <= x"0304d318";
		wait for Clk_period;
		Addr <=  "00011011100100";
		Trees_din <= x"1005e410";
		wait for Clk_period;
		Addr <=  "00011011100101";
		Trees_din <= x"15008f08";
		wait for Clk_period;
		Addr <=  "00011011100110";
		Trees_din <= x"06f67404";
		wait for Clk_period;
		Addr <=  "00011011100111";
		Trees_din <= x"00391c21";
		wait for Clk_period;
		Addr <=  "00011011101000";
		Trees_din <= x"ffbd1c21";
		wait for Clk_period;
		Addr <=  "00011011101001";
		Trees_din <= x"07005004";
		wait for Clk_period;
		Addr <=  "00011011101010";
		Trees_din <= x"00201c21";
		wait for Clk_period;
		Addr <=  "00011011101011";
		Trees_din <= x"ff8f1c21";
		wait for Clk_period;
		Addr <=  "00011011101100";
		Trees_din <= x"17016004";
		wait for Clk_period;
		Addr <=  "00011011101101";
		Trees_din <= x"fffc1c21";
		wait for Clk_period;
		Addr <=  "00011011101110";
		Trees_din <= x"00631c21";
		wait for Clk_period;
		Addr <=  "00011011101111";
		Trees_din <= x"07005910";
		wait for Clk_period;
		Addr <=  "00011011110000";
		Trees_din <= x"17039708";
		wait for Clk_period;
		Addr <=  "00011011110001";
		Trees_din <= x"1c003804";
		wait for Clk_period;
		Addr <=  "00011011110010";
		Trees_din <= x"00041c21";
		wait for Clk_period;
		Addr <=  "00011011110011";
		Trees_din <= x"ffce1c21";
		wait for Clk_period;
		Addr <=  "00011011110100";
		Trees_din <= x"0c005604";
		wait for Clk_period;
		Addr <=  "00011011110101";
		Trees_din <= x"fffe1c21";
		wait for Clk_period;
		Addr <=  "00011011110110";
		Trees_din <= x"00641c21";
		wait for Clk_period;
		Addr <=  "00011011110111";
		Trees_din <= x"00fa2408";
		wait for Clk_period;
		Addr <=  "00011011111000";
		Trees_din <= x"0f00a304";
		wait for Clk_period;
		Addr <=  "00011011111001";
		Trees_din <= x"00311c21";
		wait for Clk_period;
		Addr <=  "00011011111010";
		Trees_din <= x"ffbe1c21";
		wait for Clk_period;
		Addr <=  "00011011111011";
		Trees_din <= x"1d004404";
		wait for Clk_period;
		Addr <=  "00011011111100";
		Trees_din <= x"00001c21";
		wait for Clk_period;
		Addr <=  "00011011111101";
		Trees_din <= x"00621c21";
		wait for Clk_period;
		Addr <=  "00011011111110";
		Trees_din <= x"15009b04";
		wait for Clk_period;
		Addr <=  "00011011111111";
		Trees_din <= x"ffda1c21";
		wait for Clk_period;
		Addr <=  "00011100000000";
		Trees_din <= x"06f67804";
		wait for Clk_period;
		Addr <=  "00011100000001";
		Trees_din <= x"00131c21";
		wait for Clk_period;
		Addr <=  "00011100000010";
		Trees_din <= x"00821c21";
		wait for Clk_period;
		Addr <=  "00011100000011";
		Trees_din <= x"12035308";
		wait for Clk_period;
		Addr <=  "00011100000100";
		Trees_din <= x"0b04c104";
		wait for Clk_period;
		Addr <=  "00011100000101";
		Trees_din <= x"ff8a1c21";
		wait for Clk_period;
		Addr <=  "00011100000110";
		Trees_din <= x"ffe01c21";
		wait for Clk_period;
		Addr <=  "00011100000111";
		Trees_din <= x"00161c21";
		wait for Clk_period;
		Addr <=  "00011100001000";
		Trees_din <= x"000b1e3c";
		wait for Clk_period;
		Addr <=  "00011100001001";
		Trees_din <= x"1500b134";
		wait for Clk_period;
		Addr <=  "00011100001010";
		Trees_din <= x"20040014";
		wait for Clk_period;
		Addr <=  "00011100001011";
		Trees_din <= x"0f03fc10";
		wait for Clk_period;
		Addr <=  "00011100001100";
		Trees_din <= x"11028308";
		wait for Clk_period;
		Addr <=  "00011100001101";
		Trees_din <= x"09005804";
		wait for Clk_period;
		Addr <=  "00011100001110";
		Trees_din <= x"006a1c9d";
		wait for Clk_period;
		Addr <=  "00011100001111";
		Trees_din <= x"00061c9d";
		wait for Clk_period;
		Addr <=  "00011100010000";
		Trees_din <= x"18004204";
		wait for Clk_period;
		Addr <=  "00011100010001";
		Trees_din <= x"ffba1c9d";
		wait for Clk_period;
		Addr <=  "00011100010010";
		Trees_din <= x"00301c9d";
		wait for Clk_period;
		Addr <=  "00011100010011";
		Trees_din <= x"ffc11c9d";
		wait for Clk_period;
		Addr <=  "00011100010100";
		Trees_din <= x"0308a910";
		wait for Clk_period;
		Addr <=  "00011100010101";
		Trees_din <= x"00050808";
		wait for Clk_period;
		Addr <=  "00011100010110";
		Trees_din <= x"0800dd04";
		wait for Clk_period;
		Addr <=  "00011100010111";
		Trees_din <= x"00041c9d";
		wait for Clk_period;
		Addr <=  "00011100011000";
		Trees_din <= x"ffc41c9d";
		wait for Clk_period;
		Addr <=  "00011100011001";
		Trees_din <= x"1a00dc04";
		wait for Clk_period;
		Addr <=  "00011100011010";
		Trees_din <= x"ffeb1c9d";
		wait for Clk_period;
		Addr <=  "00011100011011";
		Trees_din <= x"005c1c9d";
		wait for Clk_period;
		Addr <=  "00011100011100";
		Trees_din <= x"08011a08";
		wait for Clk_period;
		Addr <=  "00011100011101";
		Trees_din <= x"17039104";
		wait for Clk_period;
		Addr <=  "00011100011110";
		Trees_din <= x"ffe91c9d";
		wait for Clk_period;
		Addr <=  "00011100011111";
		Trees_din <= x"00421c9d";
		wait for Clk_period;
		Addr <=  "00011100100000";
		Trees_din <= x"0e03d004";
		wait for Clk_period;
		Addr <=  "00011100100001";
		Trees_din <= x"00531c9d";
		wait for Clk_period;
		Addr <=  "00011100100010";
		Trees_din <= x"ffe01c9d";
		wait for Clk_period;
		Addr <=  "00011100100011";
		Trees_din <= x"02fdc004";
		wait for Clk_period;
		Addr <=  "00011100100100";
		Trees_din <= x"00001c9d";
		wait for Clk_period;
		Addr <=  "00011100100101";
		Trees_din <= x"ff9f1c9d";
		wait for Clk_period;
		Addr <=  "00011100100110";
		Trees_din <= x"ff961c9d";
		wait for Clk_period;
		Addr <=  "00011100100111";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00011100101000";
		Trees_din <= x"ff991d09";
		wait for Clk_period;
		Addr <=  "00011100101001";
		Trees_din <= x"1500b12c";
		wait for Clk_period;
		Addr <=  "00011100101010";
		Trees_din <= x"03075d18";
		wait for Clk_period;
		Addr <=  "00011100101011";
		Trees_din <= x"10fa2808";
		wait for Clk_period;
		Addr <=  "00011100101100";
		Trees_din <= x"08000b04";
		wait for Clk_period;
		Addr <=  "00011100101101";
		Trees_din <= x"00161d09";
		wait for Clk_period;
		Addr <=  "00011100101110";
		Trees_din <= x"ff921d09";
		wait for Clk_period;
		Addr <=  "00011100101111";
		Trees_din <= x"09005608";
		wait for Clk_period;
		Addr <=  "00011100110000";
		Trees_din <= x"1500a904";
		wait for Clk_period;
		Addr <=  "00011100110001";
		Trees_din <= x"00271d09";
		wait for Clk_period;
		Addr <=  "00011100110010";
		Trees_din <= x"ffbb1d09";
		wait for Clk_period;
		Addr <=  "00011100110011";
		Trees_din <= x"0bfb4c04";
		wait for Clk_period;
		Addr <=  "00011100110100";
		Trees_din <= x"00161d09";
		wait for Clk_period;
		Addr <=  "00011100110101";
		Trees_din <= x"ffa51d09";
		wait for Clk_period;
		Addr <=  "00011100110110";
		Trees_din <= x"16003b08";
		wait for Clk_period;
		Addr <=  "00011100110111";
		Trees_din <= x"16000104";
		wait for Clk_period;
		Addr <=  "00011100111000";
		Trees_din <= x"ffeb1d09";
		wait for Clk_period;
		Addr <=  "00011100111001";
		Trees_din <= x"00751d09";
		wait for Clk_period;
		Addr <=  "00011100111010";
		Trees_din <= x"16006d04";
		wait for Clk_period;
		Addr <=  "00011100111011";
		Trees_din <= x"ffb91d09";
		wait for Clk_period;
		Addr <=  "00011100111100";
		Trees_din <= x"0bfb1c04";
		wait for Clk_period;
		Addr <=  "00011100111101";
		Trees_din <= x"ffef1d09";
		wait for Clk_period;
		Addr <=  "00011100111110";
		Trees_din <= x"00271d09";
		wait for Clk_period;
		Addr <=  "00011100111111";
		Trees_din <= x"02fdc004";
		wait for Clk_period;
		Addr <=  "00011101000000";
		Trees_din <= x"00011d09";
		wait for Clk_period;
		Addr <=  "00011101000001";
		Trees_din <= x"ffa21d09";
		wait for Clk_period;
		Addr <=  "00011101000010";
		Trees_din <= x"0008bf2c";
		wait for Clk_period;
		Addr <=  "00011101000011";
		Trees_din <= x"0c03c424";
		wait for Clk_period;
		Addr <=  "00011101000100";
		Trees_din <= x"00063418";
		wait for Clk_period;
		Addr <=  "00011101000101";
		Trees_din <= x"0205be10";
		wait for Clk_period;
		Addr <=  "00011101000110";
		Trees_din <= x"03063408";
		wait for Clk_period;
		Addr <=  "00011101000111";
		Trees_din <= x"06f8cc04";
		wait for Clk_period;
		Addr <=  "00011101001000";
		Trees_din <= x"00061d6d";
		wait for Clk_period;
		Addr <=  "00011101001001";
		Trees_din <= x"ffa21d6d";
		wait for Clk_period;
		Addr <=  "00011101001010";
		Trees_din <= x"0c026804";
		wait for Clk_period;
		Addr <=  "00011101001011";
		Trees_din <= x"000a1d6d";
		wait for Clk_period;
		Addr <=  "00011101001100";
		Trees_din <= x"00451d6d";
		wait for Clk_period;
		Addr <=  "00011101001101";
		Trees_din <= x"16037f04";
		wait for Clk_period;
		Addr <=  "00011101001110";
		Trees_din <= x"ff961d6d";
		wait for Clk_period;
		Addr <=  "00011101001111";
		Trees_din <= x"00071d6d";
		wait for Clk_period;
		Addr <=  "00011101010000";
		Trees_din <= x"15009b04";
		wait for Clk_period;
		Addr <=  "00011101010001";
		Trees_din <= x"ffe01d6d";
		wait for Clk_period;
		Addr <=  "00011101010010";
		Trees_din <= x"1a00e304";
		wait for Clk_period;
		Addr <=  "00011101010011";
		Trees_din <= x"00741d6d";
		wait for Clk_period;
		Addr <=  "00011101010100";
		Trees_din <= x"00211d6d";
		wait for Clk_period;
		Addr <=  "00011101010101";
		Trees_din <= x"09005504";
		wait for Clk_period;
		Addr <=  "00011101010110";
		Trees_din <= x"000c1d6d";
		wait for Clk_period;
		Addr <=  "00011101010111";
		Trees_din <= x"ffa11d6d";
		wait for Clk_period;
		Addr <=  "00011101011000";
		Trees_din <= x"0f004604";
		wait for Clk_period;
		Addr <=  "00011101011001";
		Trees_din <= x"fff91d6d";
		wait for Clk_period;
		Addr <=  "00011101011010";
		Trees_din <= x"ff931d6d";
		wait for Clk_period;
		Addr <=  "00011101011011";
		Trees_din <= x"0301f914";
		wait for Clk_period;
		Addr <=  "00011101011100";
		Trees_din <= x"02031008";
		wait for Clk_period;
		Addr <=  "00011101011101";
		Trees_din <= x"10fade04";
		wait for Clk_period;
		Addr <=  "00011101011110";
		Trees_din <= x"fff41e09";
		wait for Clk_period;
		Addr <=  "00011101011111";
		Trees_din <= x"ff8e1e09";
		wait for Clk_period;
		Addr <=  "00011101100000";
		Trees_din <= x"04fd3f04";
		wait for Clk_period;
		Addr <=  "00011101100001";
		Trees_din <= x"ffad1e09";
		wait for Clk_period;
		Addr <=  "00011101100010";
		Trees_din <= x"06f52304";
		wait for Clk_period;
		Addr <=  "00011101100011";
		Trees_din <= x"ffd91e09";
		wait for Clk_period;
		Addr <=  "00011101100100";
		Trees_din <= x"00501e09";
		wait for Clk_period;
		Addr <=  "00011101100101";
		Trees_din <= x"0c002908";
		wait for Clk_period;
		Addr <=  "00011101100110";
		Trees_din <= x"1b003b04";
		wait for Clk_period;
		Addr <=  "00011101100111";
		Trees_din <= x"00031e09";
		wait for Clk_period;
		Addr <=  "00011101101000";
		Trees_din <= x"ffb01e09";
		wait for Clk_period;
		Addr <=  "00011101101001";
		Trees_din <= x"0f038420";
		wait for Clk_period;
		Addr <=  "00011101101010";
		Trees_din <= x"0f00dc10";
		wait for Clk_period;
		Addr <=  "00011101101011";
		Trees_din <= x"1900a908";
		wait for Clk_period;
		Addr <=  "00011101101100";
		Trees_din <= x"13010204";
		wait for Clk_period;
		Addr <=  "00011101101101";
		Trees_din <= x"ffef1e09";
		wait for Clk_period;
		Addr <=  "00011101101110";
		Trees_din <= x"00511e09";
		wait for Clk_period;
		Addr <=  "00011101101111";
		Trees_din <= x"06f64104";
		wait for Clk_period;
		Addr <=  "00011101110000";
		Trees_din <= x"001d1e09";
		wait for Clk_period;
		Addr <=  "00011101110001";
		Trees_din <= x"006c1e09";
		wait for Clk_period;
		Addr <=  "00011101110010";
		Trees_din <= x"11023f08";
		wait for Clk_period;
		Addr <=  "00011101110011";
		Trees_din <= x"0a015604";
		wait for Clk_period;
		Addr <=  "00011101110100";
		Trees_din <= x"00411e09";
		wait for Clk_period;
		Addr <=  "00011101110101";
		Trees_din <= x"ffe01e09";
		wait for Clk_period;
		Addr <=  "00011101110110";
		Trees_din <= x"1201f604";
		wait for Clk_period;
		Addr <=  "00011101110111";
		Trees_din <= x"00161e09";
		wait for Clk_period;
		Addr <=  "00011101111000";
		Trees_din <= x"ffa91e09";
		wait for Clk_period;
		Addr <=  "00011101111001";
		Trees_din <= x"0d002408";
		wait for Clk_period;
		Addr <=  "00011101111010";
		Trees_din <= x"06f62e04";
		wait for Clk_period;
		Addr <=  "00011101111011";
		Trees_din <= x"ffb61e09";
		wait for Clk_period;
		Addr <=  "00011101111100";
		Trees_din <= x"002c1e09";
		wait for Clk_period;
		Addr <=  "00011101111101";
		Trees_din <= x"12028708";
		wait for Clk_period;
		Addr <=  "00011101111110";
		Trees_din <= x"02fe8304";
		wait for Clk_period;
		Addr <=  "00011101111111";
		Trees_din <= x"007c1e09";
		wait for Clk_period;
		Addr <=  "00011110000000";
		Trees_din <= x"00181e09";
		wait for Clk_period;
		Addr <=  "00011110000001";
		Trees_din <= x"000b1e09";
		wait for Clk_period;
		Addr <=  "00011110000010";
		Trees_din <= x"0301f910";
		wait for Clk_period;
		Addr <=  "00011110000011";
		Trees_din <= x"07005e0c";
		wait for Clk_period;
		Addr <=  "00011110000100";
		Trees_din <= x"1b002d04";
		wait for Clk_period;
		Addr <=  "00011110000101";
		Trees_din <= x"00181ebd";
		wait for Clk_period;
		Addr <=  "00011110000110";
		Trees_din <= x"08000904";
		wait for Clk_period;
		Addr <=  "00011110000111";
		Trees_din <= x"000a1ebd";
		wait for Clk_period;
		Addr <=  "00011110001000";
		Trees_din <= x"ff851ebd";
		wait for Clk_period;
		Addr <=  "00011110001001";
		Trees_din <= x"00211ebd";
		wait for Clk_period;
		Addr <=  "00011110001010";
		Trees_din <= x"0700592c";
		wait for Clk_period;
		Addr <=  "00011110001011";
		Trees_din <= x"09005920";
		wait for Clk_period;
		Addr <=  "00011110001100";
		Trees_din <= x"08008c10";
		wait for Clk_period;
		Addr <=  "00011110001101";
		Trees_din <= x"05fa3808";
		wait for Clk_period;
		Addr <=  "00011110001110";
		Trees_din <= x"14029b04";
		wait for Clk_period;
		Addr <=  "00011110001111";
		Trees_din <= x"ffed1ebd";
		wait for Clk_period;
		Addr <=  "00011110010000";
		Trees_din <= x"005c1ebd";
		wait for Clk_period;
		Addr <=  "00011110010001";
		Trees_din <= x"07005004";
		wait for Clk_period;
		Addr <=  "00011110010010";
		Trees_din <= x"00391ebd";
		wait for Clk_period;
		Addr <=  "00011110010011";
		Trees_din <= x"ffb91ebd";
		wait for Clk_period;
		Addr <=  "00011110010100";
		Trees_din <= x"09005308";
		wait for Clk_period;
		Addr <=  "00011110010101";
		Trees_din <= x"07004a04";
		wait for Clk_period;
		Addr <=  "00011110010110";
		Trees_din <= x"00421ebd";
		wait for Clk_period;
		Addr <=  "00011110010111";
		Trees_din <= x"ffd41ebd";
		wait for Clk_period;
		Addr <=  "00011110011000";
		Trees_din <= x"0a028304";
		wait for Clk_period;
		Addr <=  "00011110011001";
		Trees_din <= x"004b1ebd";
		wait for Clk_period;
		Addr <=  "00011110011010";
		Trees_din <= x"fffa1ebd";
		wait for Clk_period;
		Addr <=  "00011110011011";
		Trees_din <= x"1a00cb08";
		wait for Clk_period;
		Addr <=  "00011110011100";
		Trees_din <= x"00feb704";
		wait for Clk_period;
		Addr <=  "00011110011101";
		Trees_din <= x"ff981ebd";
		wait for Clk_period;
		Addr <=  "00011110011110";
		Trees_din <= x"fff51ebd";
		wait for Clk_period;
		Addr <=  "00011110011111";
		Trees_din <= x"001c1ebd";
		wait for Clk_period;
		Addr <=  "00011110100000";
		Trees_din <= x"14001104";
		wait for Clk_period;
		Addr <=  "00011110100001";
		Trees_din <= x"ffcc1ebd";
		wait for Clk_period;
		Addr <=  "00011110100010";
		Trees_din <= x"1b003c10";
		wait for Clk_period;
		Addr <=  "00011110100011";
		Trees_din <= x"0306c208";
		wait for Clk_period;
		Addr <=  "00011110100100";
		Trees_din <= x"1b003704";
		wait for Clk_period;
		Addr <=  "00011110100101";
		Trees_din <= x"ffef1ebd";
		wait for Clk_period;
		Addr <=  "00011110100110";
		Trees_din <= x"ff9f1ebd";
		wait for Clk_period;
		Addr <=  "00011110100111";
		Trees_din <= x"0e02fe04";
		wait for Clk_period;
		Addr <=  "00011110101000";
		Trees_din <= x"00561ebd";
		wait for Clk_period;
		Addr <=  "00011110101001";
		Trees_din <= x"ffe11ebd";
		wait for Clk_period;
		Addr <=  "00011110101010";
		Trees_din <= x"19008908";
		wait for Clk_period;
		Addr <=  "00011110101011";
		Trees_din <= x"0200be04";
		wait for Clk_period;
		Addr <=  "00011110101100";
		Trees_din <= x"ffeb1ebd";
		wait for Clk_period;
		Addr <=  "00011110101101";
		Trees_din <= x"00401ebd";
		wait for Clk_period;
		Addr <=  "00011110101110";
		Trees_din <= x"00691ebd";
		wait for Clk_period;
		Addr <=  "00011110101111";
		Trees_din <= x"0008bf40";
		wait for Clk_period;
		Addr <=  "00011110110000";
		Trees_din <= x"00063434";
		wait for Clk_period;
		Addr <=  "00011110110001";
		Trees_din <= x"0307f520";
		wait for Clk_period;
		Addr <=  "00011110110010";
		Trees_din <= x"17000310";
		wait for Clk_period;
		Addr <=  "00011110110011";
		Trees_din <= x"1d004d08";
		wait for Clk_period;
		Addr <=  "00011110110100";
		Trees_din <= x"10045604";
		wait for Clk_period;
		Addr <=  "00011110110101";
		Trees_din <= x"ff861f49";
		wait for Clk_period;
		Addr <=  "00011110110110";
		Trees_din <= x"ffeb1f49";
		wait for Clk_period;
		Addr <=  "00011110110111";
		Trees_din <= x"20028804";
		wait for Clk_period;
		Addr <=  "00011110111000";
		Trees_din <= x"00261f49";
		wait for Clk_period;
		Addr <=  "00011110111001";
		Trees_din <= x"ffd11f49";
		wait for Clk_period;
		Addr <=  "00011110111010";
		Trees_din <= x"10052d08";
		wait for Clk_period;
		Addr <=  "00011110111011";
		Trees_din <= x"12027e04";
		wait for Clk_period;
		Addr <=  "00011110111100";
		Trees_din <= x"ffd51f49";
		wait for Clk_period;
		Addr <=  "00011110111101";
		Trees_din <= x"00261f49";
		wait for Clk_period;
		Addr <=  "00011110111110";
		Trees_din <= x"18003c04";
		wait for Clk_period;
		Addr <=  "00011110111111";
		Trees_din <= x"ffe11f49";
		wait for Clk_period;
		Addr <=  "00011111000000";
		Trees_din <= x"004e1f49";
		wait for Clk_period;
		Addr <=  "00011111000001";
		Trees_din <= x"16003b04";
		wait for Clk_period;
		Addr <=  "00011111000010";
		Trees_din <= x"00531f49";
		wait for Clk_period;
		Addr <=  "00011111000011";
		Trees_din <= x"05fde508";
		wait for Clk_period;
		Addr <=  "00011111000100";
		Trees_din <= x"05fc1204";
		wait for Clk_period;
		Addr <=  "00011111000101";
		Trees_din <= x"00011f49";
		wait for Clk_period;
		Addr <=  "00011111000110";
		Trees_din <= x"004a1f49";
		wait for Clk_period;
		Addr <=  "00011111000111";
		Trees_din <= x"0b028404";
		wait for Clk_period;
		Addr <=  "00011111001000";
		Trees_din <= x"ff911f49";
		wait for Clk_period;
		Addr <=  "00011111001001";
		Trees_din <= x"001f1f49";
		wait for Clk_period;
		Addr <=  "00011111001010";
		Trees_din <= x"15009b04";
		wait for Clk_period;
		Addr <=  "00011111001011";
		Trees_din <= x"ffe41f49";
		wait for Clk_period;
		Addr <=  "00011111001100";
		Trees_din <= x"06f77e04";
		wait for Clk_period;
		Addr <=  "00011111001101";
		Trees_din <= x"00131f49";
		wait for Clk_period;
		Addr <=  "00011111001110";
		Trees_din <= x"00691f49";
		wait for Clk_period;
		Addr <=  "00011111001111";
		Trees_din <= x"0f004604";
		wait for Clk_period;
		Addr <=  "00011111010000";
		Trees_din <= x"fffb1f49";
		wait for Clk_period;
		Addr <=  "00011111010001";
		Trees_din <= x"ff9b1f49";
		wait for Clk_period;
		Addr <=  "00011111010010";
		Trees_din <= x"03029114";
		wait for Clk_period;
		Addr <=  "00011111010011";
		Trees_din <= x"04fe3408";
		wait for Clk_period;
		Addr <=  "00011111010100";
		Trees_din <= x"04fc6e04";
		wait for Clk_period;
		Addr <=  "00011111010101";
		Trees_din <= x"ffc11fe5";
		wait for Clk_period;
		Addr <=  "00011111010110";
		Trees_din <= x"004a1fe5";
		wait for Clk_period;
		Addr <=  "00011111010111";
		Trees_din <= x"0000af08";
		wait for Clk_period;
		Addr <=  "00011111011000";
		Trees_din <= x"1d004b04";
		wait for Clk_period;
		Addr <=  "00011111011001";
		Trees_din <= x"ffc71fe5";
		wait for Clk_period;
		Addr <=  "00011111011010";
		Trees_din <= x"00331fe5";
		wait for Clk_period;
		Addr <=  "00011111011011";
		Trees_din <= x"ff8f1fe5";
		wait for Clk_period;
		Addr <=  "00011111011100";
		Trees_din <= x"09004f14";
		wait for Clk_period;
		Addr <=  "00011111011101";
		Trees_din <= x"1500b110";
		wait for Clk_period;
		Addr <=  "00011111011110";
		Trees_din <= x"0e01f00c";
		wait for Clk_period;
		Addr <=  "00011111011111";
		Trees_din <= x"0002a808";
		wait for Clk_period;
		Addr <=  "00011111100000";
		Trees_din <= x"1b003e04";
		wait for Clk_period;
		Addr <=  "00011111100001";
		Trees_din <= x"006d1fe5";
		wait for Clk_period;
		Addr <=  "00011111100010";
		Trees_din <= x"00241fe5";
		wait for Clk_period;
		Addr <=  "00011111100011";
		Trees_din <= x"000b1fe5";
		wait for Clk_period;
		Addr <=  "00011111100100";
		Trees_din <= x"fff51fe5";
		wait for Clk_period;
		Addr <=  "00011111100101";
		Trees_din <= x"ffd41fe5";
		wait for Clk_period;
		Addr <=  "00011111100110";
		Trees_din <= x"09005108";
		wait for Clk_period;
		Addr <=  "00011111100111";
		Trees_din <= x"0f008304";
		wait for Clk_period;
		Addr <=  "00011111101000";
		Trees_din <= x"00091fe5";
		wait for Clk_period;
		Addr <=  "00011111101001";
		Trees_din <= x"ffa91fe5";
		wait for Clk_period;
		Addr <=  "00011111101010";
		Trees_din <= x"01020f10";
		wait for Clk_period;
		Addr <=  "00011111101011";
		Trees_din <= x"030a7408";
		wait for Clk_period;
		Addr <=  "00011111101100";
		Trees_din <= x"00fd2504";
		wait for Clk_period;
		Addr <=  "00011111101101";
		Trees_din <= x"ffa91fe5";
		wait for Clk_period;
		Addr <=  "00011111101110";
		Trees_din <= x"fffa1fe5";
		wait for Clk_period;
		Addr <=  "00011111101111";
		Trees_din <= x"0f009a04";
		wait for Clk_period;
		Addr <=  "00011111110000";
		Trees_din <= x"ffed1fe5";
		wait for Clk_period;
		Addr <=  "00011111110001";
		Trees_din <= x"00411fe5";
		wait for Clk_period;
		Addr <=  "00011111110010";
		Trees_din <= x"06f8b808";
		wait for Clk_period;
		Addr <=  "00011111110011";
		Trees_din <= x"1201cd04";
		wait for Clk_period;
		Addr <=  "00011111110100";
		Trees_din <= x"00011fe5";
		wait for Clk_period;
		Addr <=  "00011111110101";
		Trees_din <= x"00641fe5";
		wait for Clk_period;
		Addr <=  "00011111110110";
		Trees_din <= x"02005904";
		wait for Clk_period;
		Addr <=  "00011111110111";
		Trees_din <= x"ffb91fe5";
		wait for Clk_period;
		Addr <=  "00011111111000";
		Trees_din <= x"001d1fe5";
		wait for Clk_period;
		Addr <=  "00011111111001";
		Trees_din <= x"0301f910";
		wait for Clk_period;
		Addr <=  "00011111111010";
		Trees_din <= x"07005e0c";
		wait for Clk_period;
		Addr <=  "00011111111011";
		Trees_din <= x"1b002d04";
		wait for Clk_period;
		Addr <=  "00011111111100";
		Trees_din <= x"00112071";
		wait for Clk_period;
		Addr <=  "00011111111101";
		Trees_din <= x"08000904";
		wait for Clk_period;
		Addr <=  "00011111111110";
		Trees_din <= x"00082071";
		wait for Clk_period;
		Addr <=  "00011111111111";
		Trees_din <= x"ff8c2071";
		wait for Clk_period;
		Addr <=  "00100000000000";
		Trees_din <= x"001e2071";
		wait for Clk_period;
		Addr <=  "00100000000001";
		Trees_din <= x"02053830";
		wait for Clk_period;
		Addr <=  "00100000000010";
		Trees_din <= x"0f000814";
		wait for Clk_period;
		Addr <=  "00100000000011";
		Trees_din <= x"01fc4608";
		wait for Clk_period;
		Addr <=  "00100000000100";
		Trees_din <= x"17013b04";
		wait for Clk_period;
		Addr <=  "00100000000101";
		Trees_din <= x"00492071";
		wait for Clk_period;
		Addr <=  "00100000000110";
		Trees_din <= x"fff32071";
		wait for Clk_period;
		Addr <=  "00100000000111";
		Trees_din <= x"0b004904";
		wait for Clk_period;
		Addr <=  "00100000001000";
		Trees_din <= x"00082071";
		wait for Clk_period;
		Addr <=  "00100000001001";
		Trees_din <= x"04050404";
		wait for Clk_period;
		Addr <=  "00100000001010";
		Trees_din <= x"ffe82071";
		wait for Clk_period;
		Addr <=  "00100000001011";
		Trees_din <= x"ff952071";
		wait for Clk_period;
		Addr <=  "00100000001100";
		Trees_din <= x"0f00250c";
		wait for Clk_period;
		Addr <=  "00100000001101";
		Trees_din <= x"02fd6104";
		wait for Clk_period;
		Addr <=  "00100000001110";
		Trees_din <= x"ffd92071";
		wait for Clk_period;
		Addr <=  "00100000001111";
		Trees_din <= x"15009304";
		wait for Clk_period;
		Addr <=  "00100000010000";
		Trees_din <= x"00242071";
		wait for Clk_period;
		Addr <=  "00100000010001";
		Trees_din <= x"007a2071";
		wait for Clk_period;
		Addr <=  "00100000010010";
		Trees_din <= x"0b048f08";
		wait for Clk_period;
		Addr <=  "00100000010011";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00100000010100";
		Trees_din <= x"ffce2071";
		wait for Clk_period;
		Addr <=  "00100000010101";
		Trees_din <= x"000d2071";
		wait for Clk_period;
		Addr <=  "00100000010110";
		Trees_din <= x"0b04dc04";
		wait for Clk_period;
		Addr <=  "00100000010111";
		Trees_din <= x"00672071";
		wait for Clk_period;
		Addr <=  "00100000011000";
		Trees_din <= x"00092071";
		wait for Clk_period;
		Addr <=  "00100000011001";
		Trees_din <= x"01037504";
		wait for Clk_period;
		Addr <=  "00100000011010";
		Trees_din <= x"ffa62071";
		wait for Clk_period;
		Addr <=  "00100000011011";
		Trees_din <= x"001d2071";
		wait for Clk_period;
		Addr <=  "00100000011100";
		Trees_din <= x"03075d28";
		wait for Clk_period;
		Addr <=  "00100000011101";
		Trees_din <= x"10fa2808";
		wait for Clk_period;
		Addr <=  "00100000011110";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00100000011111";
		Trees_din <= x"ff92212d";
		wait for Clk_period;
		Addr <=  "00100000100000";
		Trees_din <= x"0005212d";
		wait for Clk_period;
		Addr <=  "00100000100001";
		Trees_din <= x"0f019c10";
		wait for Clk_period;
		Addr <=  "00100000100010";
		Trees_din <= x"0108bd0c";
		wait for Clk_period;
		Addr <=  "00100000100011";
		Trees_din <= x"00fae404";
		wait for Clk_period;
		Addr <=  "00100000100100";
		Trees_din <= x"ffbb212d";
		wait for Clk_period;
		Addr <=  "00100000100101";
		Trees_din <= x"04fc6e04";
		wait for Clk_period;
		Addr <=  "00100000100110";
		Trees_din <= x"ffda212d";
		wait for Clk_period;
		Addr <=  "00100000100111";
		Trees_din <= x"0037212d";
		wait for Clk_period;
		Addr <=  "00100000101000";
		Trees_din <= x"ffa5212d";
		wait for Clk_period;
		Addr <=  "00100000101001";
		Trees_din <= x"00feee08";
		wait for Clk_period;
		Addr <=  "00100000101010";
		Trees_din <= x"00fc3a04";
		wait for Clk_period;
		Addr <=  "00100000101011";
		Trees_din <= x"ffd7212d";
		wait for Clk_period;
		Addr <=  "00100000101100";
		Trees_din <= x"004b212d";
		wait for Clk_period;
		Addr <=  "00100000101101";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00100000101110";
		Trees_din <= x"ff87212d";
		wait for Clk_period;
		Addr <=  "00100000101111";
		Trees_din <= x"0011212d";
		wait for Clk_period;
		Addr <=  "00100000110000";
		Trees_din <= x"16003b08";
		wait for Clk_period;
		Addr <=  "00100000110001";
		Trees_din <= x"06f72104";
		wait for Clk_period;
		Addr <=  "00100000110010";
		Trees_din <= x"005a212d";
		wait for Clk_period;
		Addr <=  "00100000110011";
		Trees_din <= x"0013212d";
		wait for Clk_period;
		Addr <=  "00100000110100";
		Trees_din <= x"0c015d14";
		wait for Clk_period;
		Addr <=  "00100000110101";
		Trees_din <= x"1603c908";
		wait for Clk_period;
		Addr <=  "00100000110110";
		Trees_din <= x"17002f04";
		wait for Clk_period;
		Addr <=  "00100000110111";
		Trees_din <= x"ffe9212d";
		wait for Clk_period;
		Addr <=  "00100000111000";
		Trees_din <= x"ffa2212d";
		wait for Clk_period;
		Addr <=  "00100000111001";
		Trees_din <= x"19008804";
		wait for Clk_period;
		Addr <=  "00100000111010";
		Trees_din <= x"004f212d";
		wait for Clk_period;
		Addr <=  "00100000111011";
		Trees_din <= x"05fa8c04";
		wait for Clk_period;
		Addr <=  "00100000111100";
		Trees_din <= x"002d212d";
		wait for Clk_period;
		Addr <=  "00100000111101";
		Trees_din <= x"ffde212d";
		wait for Clk_period;
		Addr <=  "00100000111110";
		Trees_din <= x"0e02100c";
		wait for Clk_period;
		Addr <=  "00100000111111";
		Trees_din <= x"01fa0f04";
		wait for Clk_period;
		Addr <=  "00100001000000";
		Trees_din <= x"ffda212d";
		wait for Clk_period;
		Addr <=  "00100001000001";
		Trees_din <= x"06f3b404";
		wait for Clk_period;
		Addr <=  "00100001000010";
		Trees_din <= x"fff5212d";
		wait for Clk_period;
		Addr <=  "00100001000011";
		Trees_din <= x"0068212d";
		wait for Clk_period;
		Addr <=  "00100001000100";
		Trees_din <= x"09005608";
		wait for Clk_period;
		Addr <=  "00100001000101";
		Trees_din <= x"08013c04";
		wait for Clk_period;
		Addr <=  "00100001000110";
		Trees_din <= x"ffb5212d";
		wait for Clk_period;
		Addr <=  "00100001000111";
		Trees_din <= x"0000212d";
		wait for Clk_period;
		Addr <=  "00100001001000";
		Trees_din <= x"00fae404";
		wait for Clk_period;
		Addr <=  "00100001001001";
		Trees_din <= x"ffe4212d";
		wait for Clk_period;
		Addr <=  "00100001001010";
		Trees_din <= x"0045212d";
		wait for Clk_period;
		Addr <=  "00100001001011";
		Trees_din <= x"0008bf38";
		wait for Clk_period;
		Addr <=  "00100001001100";
		Trees_din <= x"0c03c430";
		wait for Clk_period;
		Addr <=  "00100001001101";
		Trees_din <= x"0b04941c";
		wait for Clk_period;
		Addr <=  "00100001001110";
		Trees_din <= x"02ff0b10";
		wait for Clk_period;
		Addr <=  "00100001001111";
		Trees_din <= x"09005208";
		wait for Clk_period;
		Addr <=  "00100001010000";
		Trees_din <= x"09005004";
		wait for Clk_period;
		Addr <=  "00100001010001";
		Trees_din <= x"001321a9";
		wait for Clk_period;
		Addr <=  "00100001010010";
		Trees_din <= x"ffac21a9";
		wait for Clk_period;
		Addr <=  "00100001010011";
		Trees_din <= x"0b02fa04";
		wait for Clk_period;
		Addr <=  "00100001010100";
		Trees_din <= x"003d21a9";
		wait for Clk_period;
		Addr <=  "00100001010101";
		Trees_din <= x"fff121a9";
		wait for Clk_period;
		Addr <=  "00100001010110";
		Trees_din <= x"05ff4a08";
		wait for Clk_period;
		Addr <=  "00100001010111";
		Trees_din <= x"0c037d04";
		wait for Clk_period;
		Addr <=  "00100001011000";
		Trees_din <= x"ffd921a9";
		wait for Clk_period;
		Addr <=  "00100001011001";
		Trees_din <= x"003821a9";
		wait for Clk_period;
		Addr <=  "00100001011010";
		Trees_din <= x"003221a9";
		wait for Clk_period;
		Addr <=  "00100001011011";
		Trees_din <= x"0b04dc08";
		wait for Clk_period;
		Addr <=  "00100001011100";
		Trees_din <= x"0f003204";
		wait for Clk_period;
		Addr <=  "00100001011101";
		Trees_din <= x"ffee21a9";
		wait for Clk_period;
		Addr <=  "00100001011110";
		Trees_din <= x"006421a9";
		wait for Clk_period;
		Addr <=  "00100001011111";
		Trees_din <= x"17028008";
		wait for Clk_period;
		Addr <=  "00100001100000";
		Trees_din <= x"0d01c404";
		wait for Clk_period;
		Addr <=  "00100001100001";
		Trees_din <= x"ffe421a9";
		wait for Clk_period;
		Addr <=  "00100001100010";
		Trees_din <= x"003e21a9";
		wait for Clk_period;
		Addr <=  "00100001100011";
		Trees_din <= x"ffca21a9";
		wait for Clk_period;
		Addr <=  "00100001100100";
		Trees_din <= x"1c003304";
		wait for Clk_period;
		Addr <=  "00100001100101";
		Trees_din <= x"fff521a9";
		wait for Clk_period;
		Addr <=  "00100001100110";
		Trees_din <= x"ffb921a9";
		wait for Clk_period;
		Addr <=  "00100001100111";
		Trees_din <= x"18004204";
		wait for Clk_period;
		Addr <=  "00100001101000";
		Trees_din <= x"ffa321a9";
		wait for Clk_period;
		Addr <=  "00100001101001";
		Trees_din <= x"fffd21a9";
		wait for Clk_period;
		Addr <=  "00100001101010";
		Trees_din <= x"03075d20";
		wait for Clk_period;
		Addr <=  "00100001101011";
		Trees_din <= x"16006d08";
		wait for Clk_period;
		Addr <=  "00100001101100";
		Trees_din <= x"02ffb904";
		wait for Clk_period;
		Addr <=  "00100001101101";
		Trees_din <= x"fff3222d";
		wait for Clk_period;
		Addr <=  "00100001101110";
		Trees_din <= x"ff9b222d";
		wait for Clk_period;
		Addr <=  "00100001101111";
		Trees_din <= x"0f038414";
		wait for Clk_period;
		Addr <=  "00100001110000";
		Trees_din <= x"0f019c0c";
		wait for Clk_period;
		Addr <=  "00100001110001";
		Trees_din <= x"0108bd08";
		wait for Clk_period;
		Addr <=  "00100001110010";
		Trees_din <= x"10fa2804";
		wait for Clk_period;
		Addr <=  "00100001110011";
		Trees_din <= x"ffb6222d";
		wait for Clk_period;
		Addr <=  "00100001110100";
		Trees_din <= x"001d222d";
		wait for Clk_period;
		Addr <=  "00100001110101";
		Trees_din <= x"ffa6222d";
		wait for Clk_period;
		Addr <=  "00100001110110";
		Trees_din <= x"0efd9604";
		wait for Clk_period;
		Addr <=  "00100001110111";
		Trees_din <= x"fff6222d";
		wait for Clk_period;
		Addr <=  "00100001111000";
		Trees_din <= x"ff9b222d";
		wait for Clk_period;
		Addr <=  "00100001111001";
		Trees_din <= x"0048222d";
		wait for Clk_period;
		Addr <=  "00100001111010";
		Trees_din <= x"16003b08";
		wait for Clk_period;
		Addr <=  "00100001111011";
		Trees_din <= x"15009704";
		wait for Clk_period;
		Addr <=  "00100001111100";
		Trees_din <= x"0054222d";
		wait for Clk_period;
		Addr <=  "00100001111101";
		Trees_din <= x"000c222d";
		wait for Clk_period;
		Addr <=  "00100001111110";
		Trees_din <= x"16006d04";
		wait for Clk_period;
		Addr <=  "00100001111111";
		Trees_din <= x"ffc1222d";
		wait for Clk_period;
		Addr <=  "00100010000000";
		Trees_din <= x"19008a08";
		wait for Clk_period;
		Addr <=  "00100010000001";
		Trees_din <= x"1a00a104";
		wait for Clk_period;
		Addr <=  "00100010000010";
		Trees_din <= x"0007222d";
		wait for Clk_period;
		Addr <=  "00100010000011";
		Trees_din <= x"0059222d";
		wait for Clk_period;
		Addr <=  "00100010000100";
		Trees_din <= x"0c015d08";
		wait for Clk_period;
		Addr <=  "00100010000101";
		Trees_din <= x"0c012704";
		wait for Clk_period;
		Addr <=  "00100010000110";
		Trees_din <= x"0000222d";
		wait for Clk_period;
		Addr <=  "00100010000111";
		Trees_din <= x"ffa1222d";
		wait for Clk_period;
		Addr <=  "00100010001000";
		Trees_din <= x"1c003804";
		wait for Clk_period;
		Addr <=  "00100010001001";
		Trees_din <= x"003f222d";
		wait for Clk_period;
		Addr <=  "00100010001010";
		Trees_din <= x"ffdf222d";
		wait for Clk_period;
		Addr <=  "00100010001011";
		Trees_din <= x"03075d3c";
		wait for Clk_period;
		Addr <=  "00100010001100";
		Trees_din <= x"0101fc18";
		wait for Clk_period;
		Addr <=  "00100010001101";
		Trees_din <= x"05fd5d08";
		wait for Clk_period;
		Addr <=  "00100010001110";
		Trees_din <= x"09005104";
		wait for Clk_period;
		Addr <=  "00100010001111";
		Trees_din <= x"fff322f1";
		wait for Clk_period;
		Addr <=  "00100010010000";
		Trees_din <= x"ff9022f1";
		wait for Clk_period;
		Addr <=  "00100010010001";
		Trees_din <= x"0305c70c";
		wait for Clk_period;
		Addr <=  "00100010010010";
		Trees_din <= x"15009b04";
		wait for Clk_period;
		Addr <=  "00100010010011";
		Trees_din <= x"ffad22f1";
		wait for Clk_period;
		Addr <=  "00100010010100";
		Trees_din <= x"0800bf04";
		wait for Clk_period;
		Addr <=  "00100010010101";
		Trees_din <= x"002822f1";
		wait for Clk_period;
		Addr <=  "00100010010110";
		Trees_din <= x"fff222f1";
		wait for Clk_period;
		Addr <=  "00100010010111";
		Trees_din <= x"004322f1";
		wait for Clk_period;
		Addr <=  "00100010011000";
		Trees_din <= x"18004110";
		wait for Clk_period;
		Addr <=  "00100010011001";
		Trees_din <= x"0d01ee08";
		wait for Clk_period;
		Addr <=  "00100010011010";
		Trees_din <= x"1e006504";
		wait for Clk_period;
		Addr <=  "00100010011011";
		Trees_din <= x"ffa122f1";
		wait for Clk_period;
		Addr <=  "00100010011100";
		Trees_din <= x"fffb22f1";
		wait for Clk_period;
		Addr <=  "00100010011101";
		Trees_din <= x"1e005904";
		wait for Clk_period;
		Addr <=  "00100010011110";
		Trees_din <= x"004b22f1";
		wait for Clk_period;
		Addr <=  "00100010011111";
		Trees_din <= x"ffcd22f1";
		wait for Clk_period;
		Addr <=  "00100010100000";
		Trees_din <= x"0d02c810";
		wait for Clk_period;
		Addr <=  "00100010100001";
		Trees_din <= x"01061e08";
		wait for Clk_period;
		Addr <=  "00100010100010";
		Trees_din <= x"11009004";
		wait for Clk_period;
		Addr <=  "00100010100011";
		Trees_din <= x"001922f1";
		wait for Clk_period;
		Addr <=  "00100010100100";
		Trees_din <= x"006222f1";
		wait for Clk_period;
		Addr <=  "00100010100101";
		Trees_din <= x"0200f804";
		wait for Clk_period;
		Addr <=  "00100010100110";
		Trees_din <= x"ffd422f1";
		wait for Clk_period;
		Addr <=  "00100010100111";
		Trees_din <= x"002622f1";
		wait for Clk_period;
		Addr <=  "00100010101000";
		Trees_din <= x"ffd322f1";
		wait for Clk_period;
		Addr <=  "00100010101001";
		Trees_din <= x"0c002904";
		wait for Clk_period;
		Addr <=  "00100010101010";
		Trees_din <= x"ffcf22f1";
		wait for Clk_period;
		Addr <=  "00100010101011";
		Trees_din <= x"16003b04";
		wait for Clk_period;
		Addr <=  "00100010101100";
		Trees_din <= x"005922f1";
		wait for Clk_period;
		Addr <=  "00100010101101";
		Trees_din <= x"04041b10";
		wait for Clk_period;
		Addr <=  "00100010101110";
		Trees_din <= x"0bfb0908";
		wait for Clk_period;
		Addr <=  "00100010101111";
		Trees_din <= x"04ffc004";
		wait for Clk_period;
		Addr <=  "00100010110000";
		Trees_din <= x"002222f1";
		wait for Clk_period;
		Addr <=  "00100010110001";
		Trees_din <= x"ffce22f1";
		wait for Clk_period;
		Addr <=  "00100010110010";
		Trees_din <= x"02028904";
		wait for Clk_period;
		Addr <=  "00100010110011";
		Trees_din <= x"005222f1";
		wait for Clk_period;
		Addr <=  "00100010110100";
		Trees_din <= x"fffb22f1";
		wait for Clk_period;
		Addr <=  "00100010110101";
		Trees_din <= x"1e005e08";
		wait for Clk_period;
		Addr <=  "00100010110110";
		Trees_din <= x"0bfabb04";
		wait for Clk_period;
		Addr <=  "00100010110111";
		Trees_din <= x"ffed22f1";
		wait for Clk_period;
		Addr <=  "00100010111000";
		Trees_din <= x"005822f1";
		wait for Clk_period;
		Addr <=  "00100010111001";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00100010111010";
		Trees_din <= x"ffc722f1";
		wait for Clk_period;
		Addr <=  "00100010111011";
		Trees_din <= x"000a22f1";
		wait for Clk_period;
		Addr <=  "00100010111100";
		Trees_din <= x"030fb42c";
		wait for Clk_period;
		Addr <=  "00100010111101";
		Trees_din <= x"1500b128";
		wait for Clk_period;
		Addr <=  "00100010111110";
		Trees_din <= x"1f000220";
		wait for Clk_period;
		Addr <=  "00100010111111";
		Trees_din <= x"0304d310";
		wait for Clk_period;
		Addr <=  "00100011000000";
		Trees_din <= x"01030e08";
		wait for Clk_period;
		Addr <=  "00100011000001";
		Trees_din <= x"1603b404";
		wait for Clk_period;
		Addr <=  "00100011000010";
		Trees_din <= x"ff93234d";
		wait for Clk_period;
		Addr <=  "00100011000011";
		Trees_din <= x"ffe4234d";
		wait for Clk_period;
		Addr <=  "00100011000100";
		Trees_din <= x"0403b004";
		wait for Clk_period;
		Addr <=  "00100011000101";
		Trees_din <= x"0023234d";
		wait for Clk_period;
		Addr <=  "00100011000110";
		Trees_din <= x"ffd5234d";
		wait for Clk_period;
		Addr <=  "00100011000111";
		Trees_din <= x"06f5d408";
		wait for Clk_period;
		Addr <=  "00100011001000";
		Trees_din <= x"14018a04";
		wait for Clk_period;
		Addr <=  "00100011001001";
		Trees_din <= x"000d234d";
		wait for Clk_period;
		Addr <=  "00100011001010";
		Trees_din <= x"ffbf234d";
		wait for Clk_period;
		Addr <=  "00100011001011";
		Trees_din <= x"08022704";
		wait for Clk_period;
		Addr <=  "00100011001100";
		Trees_din <= x"0023234d";
		wait for Clk_period;
		Addr <=  "00100011001101";
		Trees_din <= x"ffd8234d";
		wait for Clk_period;
		Addr <=  "00100011001110";
		Trees_din <= x"05fafb04";
		wait for Clk_period;
		Addr <=  "00100011001111";
		Trees_din <= x"fff6234d";
		wait for Clk_period;
		Addr <=  "00100011010000";
		Trees_din <= x"0049234d";
		wait for Clk_period;
		Addr <=  "00100011010001";
		Trees_din <= x"ffc2234d";
		wait for Clk_period;
		Addr <=  "00100011010010";
		Trees_din <= x"0038234d";
		wait for Clk_period;
		Addr <=  "00100011010011";
		Trees_din <= x"0008bf38";
		wait for Clk_period;
		Addr <=  "00100011010100";
		Trees_din <= x"00063430";
		wait for Clk_period;
		Addr <=  "00100011010101";
		Trees_din <= x"00019020";
		wait for Clk_period;
		Addr <=  "00100011010110";
		Trees_din <= x"06f6d110";
		wait for Clk_period;
		Addr <=  "00100011010111";
		Trees_din <= x"0c01db08";
		wait for Clk_period;
		Addr <=  "00100011011000";
		Trees_din <= x"1b002e04";
		wait for Clk_period;
		Addr <=  "00100011011001";
		Trees_din <= x"ffe723c9";
		wait for Clk_period;
		Addr <=  "00100011011010";
		Trees_din <= x"003f23c9";
		wait for Clk_period;
		Addr <=  "00100011011011";
		Trees_din <= x"14019f04";
		wait for Clk_period;
		Addr <=  "00100011011100";
		Trees_din <= x"001f23c9";
		wait for Clk_period;
		Addr <=  "00100011011101";
		Trees_din <= x"ffc423c9";
		wait for Clk_period;
		Addr <=  "00100011011110";
		Trees_din <= x"07005308";
		wait for Clk_period;
		Addr <=  "00100011011111";
		Trees_din <= x"14011b04";
		wait for Clk_period;
		Addr <=  "00100011100000";
		Trees_din <= x"fff723c9";
		wait for Clk_period;
		Addr <=  "00100011100001";
		Trees_din <= x"004223c9";
		wait for Clk_period;
		Addr <=  "00100011100010";
		Trees_din <= x"00005104";
		wait for Clk_period;
		Addr <=  "00100011100011";
		Trees_din <= x"ffc923c9";
		wait for Clk_period;
		Addr <=  "00100011100100";
		Trees_din <= x"001e23c9";
		wait for Clk_period;
		Addr <=  "00100011100101";
		Trees_din <= x"17037c0c";
		wait for Clk_period;
		Addr <=  "00100011100110";
		Trees_din <= x"08002104";
		wait for Clk_period;
		Addr <=  "00100011100111";
		Trees_din <= x"001023c9";
		wait for Clk_period;
		Addr <=  "00100011101000";
		Trees_din <= x"0c02d404";
		wait for Clk_period;
		Addr <=  "00100011101001";
		Trees_din <= x"ff9d23c9";
		wait for Clk_period;
		Addr <=  "00100011101010";
		Trees_din <= x"fff723c9";
		wait for Clk_period;
		Addr <=  "00100011101011";
		Trees_din <= x"001e23c9";
		wait for Clk_period;
		Addr <=  "00100011101100";
		Trees_din <= x"15009b04";
		wait for Clk_period;
		Addr <=  "00100011101101";
		Trees_din <= x"ffe223c9";
		wait for Clk_period;
		Addr <=  "00100011101110";
		Trees_din <= x"004d23c9";
		wait for Clk_period;
		Addr <=  "00100011101111";
		Trees_din <= x"0f004604";
		wait for Clk_period;
		Addr <=  "00100011110000";
		Trees_din <= x"fffd23c9";
		wait for Clk_period;
		Addr <=  "00100011110001";
		Trees_din <= x"ffac23c9";
		wait for Clk_period;
		Addr <=  "00100011110010";
		Trees_din <= x"0307f534";
		wait for Clk_period;
		Addr <=  "00100011110011";
		Trees_din <= x"12fe8d10";
		wait for Clk_period;
		Addr <=  "00100011110100";
		Trees_din <= x"12fdea08";
		wait for Clk_period;
		Addr <=  "00100011110101";
		Trees_din <= x"10043004";
		wait for Clk_period;
		Addr <=  "00100011110110";
		Trees_din <= x"00112475";
		wait for Clk_period;
		Addr <=  "00100011110111";
		Trees_din <= x"ffbe2475";
		wait for Clk_period;
		Addr <=  "00100011111000";
		Trees_din <= x"12fe5804";
		wait for Clk_period;
		Addr <=  "00100011111001";
		Trees_din <= x"001c2475";
		wait for Clk_period;
		Addr <=  "00100011111010";
		Trees_din <= x"005b2475";
		wait for Clk_period;
		Addr <=  "00100011111011";
		Trees_din <= x"05ff6b20";
		wait for Clk_period;
		Addr <=  "00100011111100";
		Trees_din <= x"0e023610";
		wait for Clk_period;
		Addr <=  "00100011111101";
		Trees_din <= x"09005508";
		wait for Clk_period;
		Addr <=  "00100011111110";
		Trees_din <= x"09005404";
		wait for Clk_period;
		Addr <=  "00100011111111";
		Trees_din <= x"ffca2475";
		wait for Clk_period;
		Addr <=  "00100100000000";
		Trees_din <= x"00322475";
		wait for Clk_period;
		Addr <=  "00100100000001";
		Trees_din <= x"06f8fd04";
		wait for Clk_period;
		Addr <=  "00100100000010";
		Trees_din <= x"ff932475";
		wait for Clk_period;
		Addr <=  "00100100000011";
		Trees_din <= x"ffe42475";
		wait for Clk_period;
		Addr <=  "00100100000100";
		Trees_din <= x"09005608";
		wait for Clk_period;
		Addr <=  "00100100000101";
		Trees_din <= x"1c002b04";
		wait for Clk_period;
		Addr <=  "00100100000110";
		Trees_din <= x"00142475";
		wait for Clk_period;
		Addr <=  "00100100000111";
		Trees_din <= x"ffac2475";
		wait for Clk_period;
		Addr <=  "00100100001000";
		Trees_din <= x"07005804";
		wait for Clk_period;
		Addr <=  "00100100001001";
		Trees_din <= x"fff42475";
		wait for Clk_period;
		Addr <=  "00100100001010";
		Trees_din <= x"00432475";
		wait for Clk_period;
		Addr <=  "00100100001011";
		Trees_din <= x"00252475";
		wait for Clk_period;
		Addr <=  "00100100001100";
		Trees_din <= x"05fe1920";
		wait for Clk_period;
		Addr <=  "00100100001101";
		Trees_din <= x"0d015a0c";
		wait for Clk_period;
		Addr <=  "00100100001110";
		Trees_din <= x"1b003904";
		wait for Clk_period;
		Addr <=  "00100100001111";
		Trees_din <= x"00652475";
		wait for Clk_period;
		Addr <=  "00100100010000";
		Trees_din <= x"04041b04";
		wait for Clk_period;
		Addr <=  "00100100010001";
		Trees_din <= x"00212475";
		wait for Clk_period;
		Addr <=  "00100100010010";
		Trees_din <= x"ffde2475";
		wait for Clk_period;
		Addr <=  "00100100010011";
		Trees_din <= x"05fbcf0c";
		wait for Clk_period;
		Addr <=  "00100100010100";
		Trees_din <= x"1600e204";
		wait for Clk_period;
		Addr <=  "00100100010101";
		Trees_din <= x"00332475";
		wait for Clk_period;
		Addr <=  "00100100010110";
		Trees_din <= x"01ffd604";
		wait for Clk_period;
		Addr <=  "00100100010111";
		Trees_din <= x"ffce2475";
		wait for Clk_period;
		Addr <=  "00100100011000";
		Trees_din <= x"00132475";
		wait for Clk_period;
		Addr <=  "00100100011001";
		Trees_din <= x"01fb1904";
		wait for Clk_period;
		Addr <=  "00100100011010";
		Trees_din <= x"fff32475";
		wait for Clk_period;
		Addr <=  "00100100011011";
		Trees_din <= x"005a2475";
		wait for Clk_period;
		Addr <=  "00100100011100";
		Trees_din <= x"ffd32475";
		wait for Clk_period;
		Addr <=  "00100100011101";
		Trees_din <= x"0307f534";
		wait for Clk_period;
		Addr <=  "00100100011110";
		Trees_din <= x"12fe8d10";
		wait for Clk_period;
		Addr <=  "00100100011111";
		Trees_din <= x"12fdea08";
		wait for Clk_period;
		Addr <=  "00100100100000";
		Trees_din <= x"10043004";
		wait for Clk_period;
		Addr <=  "00100100100001";
		Trees_din <= x"00102529";
		wait for Clk_period;
		Addr <=  "00100100100010";
		Trees_din <= x"ffc32529";
		wait for Clk_period;
		Addr <=  "00100100100011";
		Trees_din <= x"12fe5804";
		wait for Clk_period;
		Addr <=  "00100100100100";
		Trees_din <= x"00192529";
		wait for Clk_period;
		Addr <=  "00100100100101";
		Trees_din <= x"00562529";
		wait for Clk_period;
		Addr <=  "00100100100110";
		Trees_din <= x"14008708";
		wait for Clk_period;
		Addr <=  "00100100100111";
		Trees_din <= x"09004e04";
		wait for Clk_period;
		Addr <=  "00100100101000";
		Trees_din <= x"00092529";
		wait for Clk_period;
		Addr <=  "00100100101001";
		Trees_din <= x"ff9c2529";
		wait for Clk_period;
		Addr <=  "00100100101010";
		Trees_din <= x"1401510c";
		wait for Clk_period;
		Addr <=  "00100100101011";
		Trees_din <= x"06f6ad04";
		wait for Clk_period;
		Addr <=  "00100100101100";
		Trees_din <= x"ffe12529";
		wait for Clk_period;
		Addr <=  "00100100101101";
		Trees_din <= x"1701ad04";
		wait for Clk_period;
		Addr <=  "00100100101110";
		Trees_din <= x"004f2529";
		wait for Clk_period;
		Addr <=  "00100100101111";
		Trees_din <= x"00062529";
		wait for Clk_period;
		Addr <=  "00100100110000";
		Trees_din <= x"01031d08";
		wait for Clk_period;
		Addr <=  "00100100110001";
		Trees_din <= x"02fea404";
		wait for Clk_period;
		Addr <=  "00100100110010";
		Trees_din <= x"fff62529";
		wait for Clk_period;
		Addr <=  "00100100110011";
		Trees_din <= x"ffa02529";
		wait for Clk_period;
		Addr <=  "00100100110100";
		Trees_din <= x"18004104";
		wait for Clk_period;
		Addr <=  "00100100110101";
		Trees_din <= x"ffd72529";
		wait for Clk_period;
		Addr <=  "00100100110110";
		Trees_din <= x"00272529";
		wait for Clk_period;
		Addr <=  "00100100110111";
		Trees_din <= x"05fe1924";
		wait for Clk_period;
		Addr <=  "00100100111000";
		Trees_din <= x"08003e08";
		wait for Clk_period;
		Addr <=  "00100100111001";
		Trees_din <= x"15009b04";
		wait for Clk_period;
		Addr <=  "00100100111010";
		Trees_din <= x"001a2529";
		wait for Clk_period;
		Addr <=  "00100100111011";
		Trees_din <= x"ffc92529";
		wait for Clk_period;
		Addr <=  "00100100111100";
		Trees_din <= x"1c00380c";
		wait for Clk_period;
		Addr <=  "00100100111101";
		Trees_din <= x"1004ee08";
		wait for Clk_period;
		Addr <=  "00100100111110";
		Trees_din <= x"11027d04";
		wait for Clk_period;
		Addr <=  "00100100111111";
		Trees_din <= x"00642529";
		wait for Clk_period;
		Addr <=  "00100101000000";
		Trees_din <= x"00212529";
		wait for Clk_period;
		Addr <=  "00100101000001";
		Trees_din <= x"fff82529";
		wait for Clk_period;
		Addr <=  "00100101000010";
		Trees_din <= x"19008908";
		wait for Clk_period;
		Addr <=  "00100101000011";
		Trees_din <= x"15008404";
		wait for Clk_period;
		Addr <=  "00100101000100";
		Trees_din <= x"fffd2529";
		wait for Clk_period;
		Addr <=  "00100101000101";
		Trees_din <= x"00402529";
		wait for Clk_period;
		Addr <=  "00100101000110";
		Trees_din <= x"05fa6e04";
		wait for Clk_period;
		Addr <=  "00100101000111";
		Trees_din <= x"00042529";
		wait for Clk_period;
		Addr <=  "00100101001000";
		Trees_din <= x"ffc72529";
		wait for Clk_period;
		Addr <=  "00100101001001";
		Trees_din <= x"ffd62529";
		wait for Clk_period;
		Addr <=  "00100101001010";
		Trees_din <= x"03029110";
		wait for Clk_period;
		Addr <=  "00100101001011";
		Trees_din <= x"04fe3408";
		wait for Clk_period;
		Addr <=  "00100101001100";
		Trees_din <= x"04fc6e04";
		wait for Clk_period;
		Addr <=  "00100101001101";
		Trees_din <= x"ffd525ad";
		wait for Clk_period;
		Addr <=  "00100101001110";
		Trees_din <= x"003825ad";
		wait for Clk_period;
		Addr <=  "00100101001111";
		Trees_din <= x"1d004c04";
		wait for Clk_period;
		Addr <=  "00100101010000";
		Trees_din <= x"ffa625ad";
		wait for Clk_period;
		Addr <=  "00100101010001";
		Trees_din <= x"000425ad";
		wait for Clk_period;
		Addr <=  "00100101010010";
		Trees_din <= x"09004c0c";
		wait for Clk_period;
		Addr <=  "00100101010011";
		Trees_din <= x"00025708";
		wait for Clk_period;
		Addr <=  "00100101010100";
		Trees_din <= x"0402ab04";
		wait for Clk_period;
		Addr <=  "00100101010101";
		Trees_din <= x"000125ad";
		wait for Clk_period;
		Addr <=  "00100101010110";
		Trees_din <= x"004d25ad";
		wait for Clk_period;
		Addr <=  "00100101010111";
		Trees_din <= x"fff425ad";
		wait for Clk_period;
		Addr <=  "00100101011000";
		Trees_din <= x"0900510c";
		wait for Clk_period;
		Addr <=  "00100101011001";
		Trees_din <= x"07005104";
		wait for Clk_period;
		Addr <=  "00100101011010";
		Trees_din <= x"001f25ad";
		wait for Clk_period;
		Addr <=  "00100101011011";
		Trees_din <= x"1201ef04";
		wait for Clk_period;
		Addr <=  "00100101011100";
		Trees_din <= x"ffef25ad";
		wait for Clk_period;
		Addr <=  "00100101011101";
		Trees_din <= x"ffaa25ad";
		wait for Clk_period;
		Addr <=  "00100101011110";
		Trees_din <= x"14007d0c";
		wait for Clk_period;
		Addr <=  "00100101011111";
		Trees_din <= x"09005708";
		wait for Clk_period;
		Addr <=  "00100101100000";
		Trees_din <= x"0308a904";
		wait for Clk_period;
		Addr <=  "00100101100001";
		Trees_din <= x"ffb525ad";
		wait for Clk_period;
		Addr <=  "00100101100010";
		Trees_din <= x"fff625ad";
		wait for Clk_period;
		Addr <=  "00100101100011";
		Trees_din <= x"001225ad";
		wait for Clk_period;
		Addr <=  "00100101100100";
		Trees_din <= x"09005708";
		wait for Clk_period;
		Addr <=  "00100101100101";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00100101100110";
		Trees_din <= x"fff025ad";
		wait for Clk_period;
		Addr <=  "00100101100111";
		Trees_din <= x"003425ad";
		wait for Clk_period;
		Addr <=  "00100101101000";
		Trees_din <= x"0e01ad04";
		wait for Clk_period;
		Addr <=  "00100101101001";
		Trees_din <= x"ffd925ad";
		wait for Clk_period;
		Addr <=  "00100101101010";
		Trees_din <= x"002325ad";
		wait for Clk_period;
		Addr <=  "00100101101011";
		Trees_din <= x"030fb434";
		wait for Clk_period;
		Addr <=  "00100101101100";
		Trees_din <= x"17039f28";
		wait for Clk_period;
		Addr <=  "00100101101101";
		Trees_din <= x"06f3bf0c";
		wait for Clk_period;
		Addr <=  "00100101101110";
		Trees_din <= x"12035308";
		wait for Clk_period;
		Addr <=  "00100101101111";
		Trees_din <= x"030a7404";
		wait for Clk_period;
		Addr <=  "00100101110000";
		Trees_din <= x"ff9e2619";
		wait for Clk_period;
		Addr <=  "00100101110001";
		Trees_din <= x"ffee2619";
		wait for Clk_period;
		Addr <=  "00100101110010";
		Trees_din <= x"00192619";
		wait for Clk_period;
		Addr <=  "00100101110011";
		Trees_din <= x"07005810";
		wait for Clk_period;
		Addr <=  "00100101110100";
		Trees_din <= x"1c003808";
		wait for Clk_period;
		Addr <=  "00100101110101";
		Trees_din <= x"12028204";
		wait for Clk_period;
		Addr <=  "00100101110110";
		Trees_din <= x"00142619";
		wait for Clk_period;
		Addr <=  "00100101110111";
		Trees_din <= x"ffca2619";
		wait for Clk_period;
		Addr <=  "00100101111000";
		Trees_din <= x"1b003f04";
		wait for Clk_period;
		Addr <=  "00100101111001";
		Trees_din <= x"ffa22619";
		wait for Clk_period;
		Addr <=  "00100101111010";
		Trees_din <= x"fff12619";
		wait for Clk_period;
		Addr <=  "00100101111011";
		Trees_din <= x"0302da04";
		wait for Clk_period;
		Addr <=  "00100101111100";
		Trees_din <= x"ffda2619";
		wait for Clk_period;
		Addr <=  "00100101111101";
		Trees_din <= x"00fcaf04";
		wait for Clk_period;
		Addr <=  "00100101111110";
		Trees_din <= x"fff12619";
		wait for Clk_period;
		Addr <=  "00100101111111";
		Trees_din <= x"00432619";
		wait for Clk_period;
		Addr <=  "00100110000000";
		Trees_din <= x"1703f108";
		wait for Clk_period;
		Addr <=  "00100110000001";
		Trees_din <= x"19009904";
		wait for Clk_period;
		Addr <=  "00100110000010";
		Trees_din <= x"00462619";
		wait for Clk_period;
		Addr <=  "00100110000011";
		Trees_din <= x"00112619";
		wait for Clk_period;
		Addr <=  "00100110000100";
		Trees_din <= x"ffd82619";
		wait for Clk_period;
		Addr <=  "00100110000101";
		Trees_din <= x"00352619";
		wait for Clk_period;
		Addr <=  "00100110000110";
		Trees_din <= x"03063420";
		wait for Clk_period;
		Addr <=  "00100110000111";
		Trees_din <= x"06fa451c";
		wait for Clk_period;
		Addr <=  "00100110001000";
		Trees_din <= x"1500a918";
		wait for Clk_period;
		Addr <=  "00100110001001";
		Trees_din <= x"0403780c";
		wait for Clk_period;
		Addr <=  "00100110001010";
		Trees_din <= x"09005708";
		wait for Clk_period;
		Addr <=  "00100110001011";
		Trees_din <= x"01029904";
		wait for Clk_period;
		Addr <=  "00100110001100";
		Trees_din <= x"fff226a5";
		wait for Clk_period;
		Addr <=  "00100110001101";
		Trees_din <= x"004826a5";
		wait for Clk_period;
		Addr <=  "00100110001110";
		Trees_din <= x"ffe126a5";
		wait for Clk_period;
		Addr <=  "00100110001111";
		Trees_din <= x"10054a08";
		wait for Clk_period;
		Addr <=  "00100110010000";
		Trees_din <= x"06f6ad04";
		wait for Clk_period;
		Addr <=  "00100110010001";
		Trees_din <= x"ffbb26a5";
		wait for Clk_period;
		Addr <=  "00100110010010";
		Trees_din <= x"000e26a5";
		wait for Clk_period;
		Addr <=  "00100110010011";
		Trees_din <= x"002326a5";
		wait for Clk_period;
		Addr <=  "00100110010100";
		Trees_din <= x"ffae26a5";
		wait for Clk_period;
		Addr <=  "00100110010101";
		Trees_din <= x"ffb326a5";
		wait for Clk_period;
		Addr <=  "00100110010110";
		Trees_din <= x"15008208";
		wait for Clk_period;
		Addr <=  "00100110010111";
		Trees_din <= x"1100e804";
		wait for Clk_period;
		Addr <=  "00100110011000";
		Trees_din <= x"ffc326a5";
		wait for Clk_period;
		Addr <=  "00100110011001";
		Trees_din <= x"000126a5";
		wait for Clk_period;
		Addr <=  "00100110011010";
		Trees_din <= x"19008904";
		wait for Clk_period;
		Addr <=  "00100110011011";
		Trees_din <= x"004726a5";
		wait for Clk_period;
		Addr <=  "00100110011100";
		Trees_din <= x"1100fa0c";
		wait for Clk_period;
		Addr <=  "00100110011101";
		Trees_din <= x"07005608";
		wait for Clk_period;
		Addr <=  "00100110011110";
		Trees_din <= x"06f7b304";
		wait for Clk_period;
		Addr <=  "00100110011111";
		Trees_din <= x"ffd526a5";
		wait for Clk_period;
		Addr <=  "00100110100000";
		Trees_din <= x"004326a5";
		wait for Clk_period;
		Addr <=  "00100110100001";
		Trees_din <= x"004f26a5";
		wait for Clk_period;
		Addr <=  "00100110100010";
		Trees_din <= x"1b002f08";
		wait for Clk_period;
		Addr <=  "00100110100011";
		Trees_din <= x"0bfa8104";
		wait for Clk_period;
		Addr <=  "00100110100100";
		Trees_din <= x"ffe226a5";
		wait for Clk_period;
		Addr <=  "00100110100101";
		Trees_din <= x"004926a5";
		wait for Clk_period;
		Addr <=  "00100110100110";
		Trees_din <= x"01fa9904";
		wait for Clk_period;
		Addr <=  "00100110100111";
		Trees_din <= x"002026a5";
		wait for Clk_period;
		Addr <=  "00100110101000";
		Trees_din <= x"ffe126a5";
		wait for Clk_period;
		Addr <=  "00100110101001";
		Trees_din <= x"0307f534";
		wait for Clk_period;
		Addr <=  "00100110101010";
		Trees_din <= x"12fe8d10";
		wait for Clk_period;
		Addr <=  "00100110101011";
		Trees_din <= x"12fdea08";
		wait for Clk_period;
		Addr <=  "00100110101100";
		Trees_din <= x"02ff2a04";
		wait for Clk_period;
		Addr <=  "00100110101101";
		Trees_din <= x"000f2751";
		wait for Clk_period;
		Addr <=  "00100110101110";
		Trees_din <= x"ffce2751";
		wait for Clk_period;
		Addr <=  "00100110101111";
		Trees_din <= x"12fe5804";
		wait for Clk_period;
		Addr <=  "00100110110000";
		Trees_din <= x"00122751";
		wait for Clk_period;
		Addr <=  "00100110110001";
		Trees_din <= x"004c2751";
		wait for Clk_period;
		Addr <=  "00100110110010";
		Trees_din <= x"05ff4a20";
		wait for Clk_period;
		Addr <=  "00100110110011";
		Trees_din <= x"0e023610";
		wait for Clk_period;
		Addr <=  "00100110110100";
		Trees_din <= x"1900a108";
		wait for Clk_period;
		Addr <=  "00100110110101";
		Trees_din <= x"1500a104";
		wait for Clk_period;
		Addr <=  "00100110110110";
		Trees_din <= x"ffac2751";
		wait for Clk_period;
		Addr <=  "00100110110111";
		Trees_din <= x"00062751";
		wait for Clk_period;
		Addr <=  "00100110111000";
		Trees_din <= x"0effcc04";
		wait for Clk_period;
		Addr <=  "00100110111001";
		Trees_din <= x"00322751";
		wait for Clk_period;
		Addr <=  "00100110111010";
		Trees_din <= x"ffc22751";
		wait for Clk_period;
		Addr <=  "00100110111011";
		Trees_din <= x"05fbb608";
		wait for Clk_period;
		Addr <=  "00100110111100";
		Trees_din <= x"10fb0104";
		wait for Clk_period;
		Addr <=  "00100110111101";
		Trees_din <= x"003b2751";
		wait for Clk_period;
		Addr <=  "00100110111110";
		Trees_din <= x"fff82751";
		wait for Clk_period;
		Addr <=  "00100110111111";
		Trees_din <= x"06f71604";
		wait for Clk_period;
		Addr <=  "00100111000000";
		Trees_din <= x"ffb02751";
		wait for Clk_period;
		Addr <=  "00100111000001";
		Trees_din <= x"00102751";
		wait for Clk_period;
		Addr <=  "00100111000010";
		Trees_din <= x"001d2751";
		wait for Clk_period;
		Addr <=  "00100111000011";
		Trees_din <= x"05fde520";
		wait for Clk_period;
		Addr <=  "00100111000100";
		Trees_din <= x"08003e08";
		wait for Clk_period;
		Addr <=  "00100111000101";
		Trees_din <= x"15009b04";
		wait for Clk_period;
		Addr <=  "00100111000110";
		Trees_din <= x"00172751";
		wait for Clk_period;
		Addr <=  "00100111000111";
		Trees_din <= x"ffce2751";
		wait for Clk_period;
		Addr <=  "00100111001000";
		Trees_din <= x"1c00380c";
		wait for Clk_period;
		Addr <=  "00100111001001";
		Trees_din <= x"13fa6404";
		wait for Clk_period;
		Addr <=  "00100111001010";
		Trees_din <= x"fffc2751";
		wait for Clk_period;
		Addr <=  "00100111001011";
		Trees_din <= x"0e021004";
		wait for Clk_period;
		Addr <=  "00100111001100";
		Trees_din <= x"00662751";
		wait for Clk_period;
		Addr <=  "00100111001101";
		Trees_din <= x"001e2751";
		wait for Clk_period;
		Addr <=  "00100111001110";
		Trees_din <= x"030a7404";
		wait for Clk_period;
		Addr <=  "00100111001111";
		Trees_din <= x"ffd02751";
		wait for Clk_period;
		Addr <=  "00100111010000";
		Trees_din <= x"13ffeb04";
		wait for Clk_period;
		Addr <=  "00100111010001";
		Trees_din <= x"003b2751";
		wait for Clk_period;
		Addr <=  "00100111010010";
		Trees_din <= x"ffe82751";
		wait for Clk_period;
		Addr <=  "00100111010011";
		Trees_din <= x"ffde2751";
		wait for Clk_period;
		Addr <=  "00100111010100";
		Trees_din <= x"03029110";
		wait for Clk_period;
		Addr <=  "00100111010101";
		Trees_din <= x"04fe3408";
		wait for Clk_period;
		Addr <=  "00100111010110";
		Trees_din <= x"04fc6e04";
		wait for Clk_period;
		Addr <=  "00100111010111";
		Trees_din <= x"ffd727cd";
		wait for Clk_period;
		Addr <=  "00100111011000";
		Trees_din <= x"002f27cd";
		wait for Clk_period;
		Addr <=  "00100111011001";
		Trees_din <= x"0000af04";
		wait for Clk_period;
		Addr <=  "00100111011010";
		Trees_din <= x"000027cd";
		wait for Clk_period;
		Addr <=  "00100111011011";
		Trees_din <= x"ffa627cd";
		wait for Clk_period;
		Addr <=  "00100111011100";
		Trees_din <= x"0205382c";
		wait for Clk_period;
		Addr <=  "00100111011101";
		Trees_din <= x"0f00090c";
		wait for Clk_period;
		Addr <=  "00100111011110";
		Trees_din <= x"01fc4604";
		wait for Clk_period;
		Addr <=  "00100111011111";
		Trees_din <= x"001627cd";
		wait for Clk_period;
		Addr <=  "00100111100000";
		Trees_din <= x"0b004904";
		wait for Clk_period;
		Addr <=  "00100111100001";
		Trees_din <= x"000d27cd";
		wait for Clk_period;
		Addr <=  "00100111100010";
		Trees_din <= x"ffb727cd";
		wait for Clk_period;
		Addr <=  "00100111100011";
		Trees_din <= x"0f00dc10";
		wait for Clk_period;
		Addr <=  "00100111100100";
		Trees_din <= x"02fdc008";
		wait for Clk_period;
		Addr <=  "00100111100101";
		Trees_din <= x"0b03a104";
		wait for Clk_period;
		Addr <=  "00100111100110";
		Trees_din <= x"002527cd";
		wait for Clk_period;
		Addr <=  "00100111100111";
		Trees_din <= x"ffd627cd";
		wait for Clk_period;
		Addr <=  "00100111101000";
		Trees_din <= x"0bf9ce04";
		wait for Clk_period;
		Addr <=  "00100111101001";
		Trees_din <= x"fffc27cd";
		wait for Clk_period;
		Addr <=  "00100111101010";
		Trees_din <= x"004427cd";
		wait for Clk_period;
		Addr <=  "00100111101011";
		Trees_din <= x"02002408";
		wait for Clk_period;
		Addr <=  "00100111101100";
		Trees_din <= x"14015804";
		wait for Clk_period;
		Addr <=  "00100111101101";
		Trees_din <= x"ffce27cd";
		wait for Clk_period;
		Addr <=  "00100111101110";
		Trees_din <= x"002a27cd";
		wait for Clk_period;
		Addr <=  "00100111101111";
		Trees_din <= x"0d030504";
		wait for Clk_period;
		Addr <=  "00100111110000";
		Trees_din <= x"ffb327cd";
		wait for Clk_period;
		Addr <=  "00100111110001";
		Trees_din <= x"003827cd";
		wait for Clk_period;
		Addr <=  "00100111110010";
		Trees_din <= x"ffd027cd";
		wait for Clk_period;
		Addr <=  "00100111110011";
		Trees_din <= x"03063420";
		wait for Clk_period;
		Addr <=  "00100111110100";
		Trees_din <= x"1500a91c";
		wait for Clk_period;
		Addr <=  "00100111110101";
		Trees_din <= x"06fa4518";
		wait for Clk_period;
		Addr <=  "00100111110110";
		Trees_din <= x"0f019c0c";
		wait for Clk_period;
		Addr <=  "00100111110111";
		Trees_din <= x"1c003d08";
		wait for Clk_period;
		Addr <=  "00100111111000";
		Trees_din <= x"0105d004";
		wait for Clk_period;
		Addr <=  "00100111111001";
		Trees_din <= x"00382849";
		wait for Clk_period;
		Addr <=  "00100111111010";
		Trees_din <= x"fff62849";
		wait for Clk_period;
		Addr <=  "00100111111011";
		Trees_din <= x"ffda2849";
		wait for Clk_period;
		Addr <=  "00100111111100";
		Trees_din <= x"05fac804";
		wait for Clk_period;
		Addr <=  "00100111111101";
		Trees_din <= x"00242849";
		wait for Clk_period;
		Addr <=  "00100111111110";
		Trees_din <= x"16007004";
		wait for Clk_period;
		Addr <=  "00100111111111";
		Trees_din <= x"ffe92849";
		wait for Clk_period;
		Addr <=  "00101000000000";
		Trees_din <= x"ffa82849";
		wait for Clk_period;
		Addr <=  "00101000000001";
		Trees_din <= x"ffbc2849";
		wait for Clk_period;
		Addr <=  "00101000000010";
		Trees_din <= x"ffb42849";
		wait for Clk_period;
		Addr <=  "00101000000011";
		Trees_din <= x"15008208";
		wait for Clk_period;
		Addr <=  "00101000000100";
		Trees_din <= x"17007904";
		wait for Clk_period;
		Addr <=  "00101000000101";
		Trees_din <= x"ffca2849";
		wait for Clk_period;
		Addr <=  "00101000000110";
		Trees_din <= x"00002849";
		wait for Clk_period;
		Addr <=  "00101000000111";
		Trees_din <= x"15009008";
		wait for Clk_period;
		Addr <=  "00101000001000";
		Trees_din <= x"02010804";
		wait for Clk_period;
		Addr <=  "00101000001001";
		Trees_din <= x"005c2849";
		wait for Clk_period;
		Addr <=  "00101000001010";
		Trees_din <= x"ffde2849";
		wait for Clk_period;
		Addr <=  "00101000001011";
		Trees_din <= x"15009504";
		wait for Clk_period;
		Addr <=  "00101000001100";
		Trees_din <= x"ffce2849";
		wait for Clk_period;
		Addr <=  "00101000001101";
		Trees_din <= x"08003e04";
		wait for Clk_period;
		Addr <=  "00101000001110";
		Trees_din <= x"ffe62849";
		wait for Clk_period;
		Addr <=  "00101000001111";
		Trees_din <= x"19009704";
		wait for Clk_period;
		Addr <=  "00101000010000";
		Trees_din <= x"004e2849";
		wait for Clk_period;
		Addr <=  "00101000010001";
		Trees_din <= x"000f2849";
		wait for Clk_period;
		Addr <=  "00101000010010";
		Trees_din <= x"0008bf4c";
		wait for Clk_period;
		Addr <=  "00101000010011";
		Trees_din <= x"04025d20";
		wait for Clk_period;
		Addr <=  "00101000010100";
		Trees_din <= x"02fe7808";
		wait for Clk_period;
		Addr <=  "00101000010101";
		Trees_din <= x"16032104";
		wait for Clk_period;
		Addr <=  "00101000010110";
		Trees_din <= x"000d28e5";
		wait for Clk_period;
		Addr <=  "00101000010111";
		Trees_din <= x"ffcf28e5";
		wait for Clk_period;
		Addr <=  "00101000011000";
		Trees_din <= x"13ffcd10";
		wait for Clk_period;
		Addr <=  "00101000011001";
		Trees_din <= x"02031e08";
		wait for Clk_period;
		Addr <=  "00101000011010";
		Trees_din <= x"1004e304";
		wait for Clk_period;
		Addr <=  "00101000011011";
		Trees_din <= x"005428e5";
		wait for Clk_period;
		Addr <=  "00101000011100";
		Trees_din <= x"001328e5";
		wait for Clk_period;
		Addr <=  "00101000011101";
		Trees_din <= x"11000d04";
		wait for Clk_period;
		Addr <=  "00101000011110";
		Trees_din <= x"003f28e5";
		wait for Clk_period;
		Addr <=  "00101000011111";
		Trees_din <= x"ffe128e5";
		wait for Clk_period;
		Addr <=  "00101000100000";
		Trees_din <= x"00011804";
		wait for Clk_period;
		Addr <=  "00101000100001";
		Trees_din <= x"001428e5";
		wait for Clk_period;
		Addr <=  "00101000100010";
		Trees_din <= x"ffd728e5";
		wait for Clk_period;
		Addr <=  "00101000100011";
		Trees_din <= x"02fe6214";
		wait for Clk_period;
		Addr <=  "00101000100100";
		Trees_din <= x"17000008";
		wait for Clk_period;
		Addr <=  "00101000100101";
		Trees_din <= x"16003904";
		wait for Clk_period;
		Addr <=  "00101000100110";
		Trees_din <= x"002028e5";
		wait for Clk_period;
		Addr <=  "00101000100111";
		Trees_din <= x"ffab28e5";
		wait for Clk_period;
		Addr <=  "00101000101000";
		Trees_din <= x"13fa6404";
		wait for Clk_period;
		Addr <=  "00101000101001";
		Trees_din <= x"fff128e5";
		wait for Clk_period;
		Addr <=  "00101000101010";
		Trees_din <= x"0d030104";
		wait for Clk_period;
		Addr <=  "00101000101011";
		Trees_din <= x"004d28e5";
		wait for Clk_period;
		Addr <=  "00101000101100";
		Trees_din <= x"fffa28e5";
		wait for Clk_period;
		Addr <=  "00101000101101";
		Trees_din <= x"00001410";
		wait for Clk_period;
		Addr <=  "00101000101110";
		Trees_din <= x"00fc3a08";
		wait for Clk_period;
		Addr <=  "00101000101111";
		Trees_din <= x"030a7404";
		wait for Clk_period;
		Addr <=  "00101000110000";
		Trees_din <= x"ffc228e5";
		wait for Clk_period;
		Addr <=  "00101000110001";
		Trees_din <= x"001028e5";
		wait for Clk_period;
		Addr <=  "00101000110010";
		Trees_din <= x"19009f04";
		wait for Clk_period;
		Addr <=  "00101000110011";
		Trees_din <= x"004128e5";
		wait for Clk_period;
		Addr <=  "00101000110100";
		Trees_din <= x"ffe028e5";
		wait for Clk_period;
		Addr <=  "00101000110101";
		Trees_din <= x"0d027a04";
		wait for Clk_period;
		Addr <=  "00101000110110";
		Trees_din <= x"ffa928e5";
		wait for Clk_period;
		Addr <=  "00101000110111";
		Trees_din <= x"fff128e5";
		wait for Clk_period;
		Addr <=  "00101000111000";
		Trees_din <= x"ffcf28e5";
		wait for Clk_period;
		Addr <=  "00101000111001";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  3
        -----------
		Addr <=  "00000000000000";
		Trees_din <= x"0406be3c";
		wait for Clk_period;
		Addr <=  "00000000000001";
		Trees_din <= x"04045e20";
		wait for Clk_period;
		Addr <=  "00000000000010";
		Trees_din <= x"0401dd04";
		wait for Clk_period;
		Addr <=  "00000000000011";
		Trees_din <= x"ff4f0125";
		wait for Clk_period;
		Addr <=  "00000000000100";
		Trees_din <= x"0efcb00c";
		wait for Clk_period;
		Addr <=  "00000000000101";
		Trees_din <= x"17005708";
		wait for Clk_period;
		Addr <=  "00000000000110";
		Trees_din <= x"18004804";
		wait for Clk_period;
		Addr <=  "00000000000111";
		Trees_din <= x"ff640125";
		wait for Clk_period;
		Addr <=  "00000000001000";
		Trees_din <= x"00590125";
		wait for Clk_period;
		Addr <=  "00000000001001";
		Trees_din <= x"013c0125";
		wait for Clk_period;
		Addr <=  "00000000001010";
		Trees_din <= x"04025d08";
		wait for Clk_period;
		Addr <=  "00000000001011";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00000000001100";
		Trees_din <= x"006b0125";
		wait for Clk_period;
		Addr <=  "00000000001101";
		Trees_din <= x"ff7d0125";
		wait for Clk_period;
		Addr <=  "00000000001110";
		Trees_din <= x"05feb404";
		wait for Clk_period;
		Addr <=  "00000000001111";
		Trees_din <= x"ff500125";
		wait for Clk_period;
		Addr <=  "00000000010000";
		Trees_din <= x"ffa70125";
		wait for Clk_period;
		Addr <=  "00000000010001";
		Trees_din <= x"0c03f818";
		wait for Clk_period;
		Addr <=  "00000000010010";
		Trees_din <= x"11046110";
		wait for Clk_period;
		Addr <=  "00000000010011";
		Trees_din <= x"06f55708";
		wait for Clk_period;
		Addr <=  "00000000010100";
		Trees_din <= x"12ffbe04";
		wait for Clk_period;
		Addr <=  "00000000010101";
		Trees_din <= x"ffc00125";
		wait for Clk_period;
		Addr <=  "00000000010110";
		Trees_din <= x"ff560125";
		wait for Clk_period;
		Addr <=  "00000000010111";
		Trees_din <= x"1c003404";
		wait for Clk_period;
		Addr <=  "00000000011000";
		Trees_din <= x"008e0125";
		wait for Clk_period;
		Addr <=  "00000000011001";
		Trees_din <= x"ff9d0125";
		wait for Clk_period;
		Addr <=  "00000000011010";
		Trees_din <= x"05fbe604";
		wait for Clk_period;
		Addr <=  "00000000011011";
		Trees_din <= x"fff10125";
		wait for Clk_period;
		Addr <=  "00000000011100";
		Trees_din <= x"02500125";
		wait for Clk_period;
		Addr <=  "00000000011101";
		Trees_din <= x"01c50125";
		wait for Clk_period;
		Addr <=  "00000000011110";
		Trees_din <= x"040a4a38";
		wait for Clk_period;
		Addr <=  "00000000011111";
		Trees_din <= x"05fcf120";
		wait for Clk_period;
		Addr <=  "00000000100000";
		Trees_din <= x"030a7410";
		wait for Clk_period;
		Addr <=  "00000000100001";
		Trees_din <= x"03fd0608";
		wait for Clk_period;
		Addr <=  "00000000100010";
		Trees_din <= x"00fd2504";
		wait for Clk_period;
		Addr <=  "00000000100011";
		Trees_din <= x"00270125";
		wait for Clk_period;
		Addr <=  "00000000100100";
		Trees_din <= x"ff6e0125";
		wait for Clk_period;
		Addr <=  "00000000100101";
		Trees_din <= x"15007b04";
		wait for Clk_period;
		Addr <=  "00000000100110";
		Trees_din <= x"ff7a0125";
		wait for Clk_period;
		Addr <=  "00000000100111";
		Trees_din <= x"01290125";
		wait for Clk_period;
		Addr <=  "00000000101000";
		Trees_din <= x"13004e08";
		wait for Clk_period;
		Addr <=  "00000000101001";
		Trees_din <= x"08005104";
		wait for Clk_period;
		Addr <=  "00000000101010";
		Trees_din <= x"00270125";
		wait for Clk_period;
		Addr <=  "00000000101011";
		Trees_din <= x"ff5f0125";
		wait for Clk_period;
		Addr <=  "00000000101100";
		Trees_din <= x"14010404";
		wait for Clk_period;
		Addr <=  "00000000101101";
		Trees_din <= x"ff9d0125";
		wait for Clk_period;
		Addr <=  "00000000101110";
		Trees_din <= x"013c0125";
		wait for Clk_period;
		Addr <=  "00000000101111";
		Trees_din <= x"18004a10";
		wait for Clk_period;
		Addr <=  "00000000110000";
		Trees_din <= x"01fdac08";
		wait for Clk_period;
		Addr <=  "00000000110001";
		Trees_din <= x"1101b604";
		wait for Clk_period;
		Addr <=  "00000000110010";
		Trees_din <= x"ff890125";
		wait for Clk_period;
		Addr <=  "00000000110011";
		Trees_din <= x"01f80125";
		wait for Clk_period;
		Addr <=  "00000000110100";
		Trees_din <= x"01038904";
		wait for Clk_period;
		Addr <=  "00000000110101";
		Trees_din <= x"02fa0125";
		wait for Clk_period;
		Addr <=  "00000000110110";
		Trees_din <= x"00b20125";
		wait for Clk_period;
		Addr <=  "00000000110111";
		Trees_din <= x"1100b304";
		wait for Clk_period;
		Addr <=  "00000000111000";
		Trees_din <= x"013c0125";
		wait for Clk_period;
		Addr <=  "00000000111001";
		Trees_din <= x"ff850125";
		wait for Clk_period;
		Addr <=  "00000000111010";
		Trees_din <= x"030a7418";
		wait for Clk_period;
		Addr <=  "00000000111011";
		Trees_din <= x"0202d90c";
		wait for Clk_period;
		Addr <=  "00000000111100";
		Trees_din <= x"010a4208";
		wait for Clk_period;
		Addr <=  "00000000111101";
		Trees_din <= x"040b2e04";
		wait for Clk_period;
		Addr <=  "00000000111110";
		Trees_din <= x"01f40125";
		wait for Clk_period;
		Addr <=  "00000000111111";
		Trees_din <= x"03a30125";
		wait for Clk_period;
		Addr <=  "00000001000000";
		Trees_din <= x"00c10125";
		wait for Clk_period;
		Addr <=  "00000001000001";
		Trees_din <= x"11019508";
		wait for Clk_period;
		Addr <=  "00000001000010";
		Trees_din <= x"0a02a204";
		wait for Clk_period;
		Addr <=  "00000001000011";
		Trees_din <= x"02600125";
		wait for Clk_period;
		Addr <=  "00000001000100";
		Trees_din <= x"00120125";
		wait for Clk_period;
		Addr <=  "00000001000101";
		Trees_din <= x"ff950125";
		wait for Clk_period;
		Addr <=  "00000001000110";
		Trees_din <= x"0b02fa04";
		wait for Clk_period;
		Addr <=  "00000001000111";
		Trees_din <= x"ff6c0125";
		wait for Clk_period;
		Addr <=  "00000001001000";
		Trees_din <= x"01290125";
		wait for Clk_period;
		Addr <=  "00000001001001";
		Trees_din <= x"0406be54";
		wait for Clk_period;
		Addr <=  "00000001001010";
		Trees_din <= x"04041b2c";
		wait for Clk_period;
		Addr <=  "00000001001011";
		Trees_din <= x"0401dd10";
		wait for Clk_period;
		Addr <=  "00000001001100";
		Trees_din <= x"03fbf604";
		wait for Clk_period;
		Addr <=  "00000001001101";
		Trees_din <= x"ff540249";
		wait for Clk_period;
		Addr <=  "00000001001110";
		Trees_din <= x"0f040008";
		wait for Clk_period;
		Addr <=  "00000001001111";
		Trees_din <= x"0e045b04";
		wait for Clk_period;
		Addr <=  "00000001010000";
		Trees_din <= x"ff5c0249";
		wait for Clk_period;
		Addr <=  "00000001010001";
		Trees_din <= x"ffc70249";
		wait for Clk_period;
		Addr <=  "00000001010010";
		Trees_din <= x"00410249";
		wait for Clk_period;
		Addr <=  "00000001010011";
		Trees_din <= x"05fd7a0c";
		wait for Clk_period;
		Addr <=  "00000001010100";
		Trees_din <= x"13f85404";
		wait for Clk_period;
		Addr <=  "00000001010101";
		Trees_din <= x"00240249";
		wait for Clk_period;
		Addr <=  "00000001010110";
		Trees_din <= x"1a008d04";
		wait for Clk_period;
		Addr <=  "00000001010111";
		Trees_din <= x"000b0249";
		wait for Clk_period;
		Addr <=  "00000001011000";
		Trees_din <= x"ff5d0249";
		wait for Clk_period;
		Addr <=  "00000001011001";
		Trees_din <= x"15009c08";
		wait for Clk_period;
		Addr <=  "00000001011010";
		Trees_din <= x"03fcb704";
		wait for Clk_period;
		Addr <=  "00000001011011";
		Trees_din <= x"00230249";
		wait for Clk_period;
		Addr <=  "00000001011100";
		Trees_din <= x"ff620249";
		wait for Clk_period;
		Addr <=  "00000001011101";
		Trees_din <= x"0d024404";
		wait for Clk_period;
		Addr <=  "00000001011110";
		Trees_din <= x"ff870249";
		wait for Clk_period;
		Addr <=  "00000001011111";
		Trees_din <= x"014b0249";
		wait for Clk_period;
		Addr <=  "00000001100000";
		Trees_din <= x"06f4ea10";
		wait for Clk_period;
		Addr <=  "00000001100001";
		Trees_din <= x"1104610c";
		wait for Clk_period;
		Addr <=  "00000001100010";
		Trees_din <= x"12ffbe08";
		wait for Clk_period;
		Addr <=  "00000001100011";
		Trees_din <= x"0afda204";
		wait for Clk_period;
		Addr <=  "00000001100100";
		Trees_din <= x"00cb0249";
		wait for Clk_period;
		Addr <=  "00000001100101";
		Trees_din <= x"ff6d0249";
		wait for Clk_period;
		Addr <=  "00000001100110";
		Trees_din <= x"ff5d0249";
		wait for Clk_period;
		Addr <=  "00000001100111";
		Trees_din <= x"00a20249";
		wait for Clk_period;
		Addr <=  "00000001101000";
		Trees_din <= x"0308a910";
		wait for Clk_period;
		Addr <=  "00000001101001";
		Trees_din <= x"0c024e08";
		wait for Clk_period;
		Addr <=  "00000001101010";
		Trees_din <= x"1e006404";
		wait for Clk_period;
		Addr <=  "00000001101011";
		Trees_din <= x"009e0249";
		wait for Clk_period;
		Addr <=  "00000001101100";
		Trees_din <= x"ff890249";
		wait for Clk_period;
		Addr <=  "00000001101101";
		Trees_din <= x"12007b04";
		wait for Clk_period;
		Addr <=  "00000001101110";
		Trees_din <= x"ff8e0249";
		wait for Clk_period;
		Addr <=  "00000001101111";
		Trees_din <= x"01a00249";
		wait for Clk_period;
		Addr <=  "00000001110000";
		Trees_din <= x"10050404";
		wait for Clk_period;
		Addr <=  "00000001110001";
		Trees_din <= x"ff600249";
		wait for Clk_period;
		Addr <=  "00000001110010";
		Trees_din <= x"00560249";
		wait for Clk_period;
		Addr <=  "00000001110011";
		Trees_din <= x"030a7428";
		wait for Clk_period;
		Addr <=  "00000001110100";
		Trees_din <= x"0205511c";
		wait for Clk_period;
		Addr <=  "00000001110101";
		Trees_din <= x"01084110";
		wait for Clk_period;
		Addr <=  "00000001110110";
		Trees_din <= x"18004208";
		wait for Clk_period;
		Addr <=  "00000001110111";
		Trees_din <= x"07004804";
		wait for Clk_period;
		Addr <=  "00000001111000";
		Trees_din <= x"002c0249";
		wait for Clk_period;
		Addr <=  "00000001111001";
		Trees_din <= x"01a90249";
		wait for Clk_period;
		Addr <=  "00000001111010";
		Trees_din <= x"05fbd904";
		wait for Clk_period;
		Addr <=  "00000001111011";
		Trees_din <= x"017e0249";
		wait for Clk_period;
		Addr <=  "00000001111100";
		Trees_din <= x"00a00249";
		wait for Clk_period;
		Addr <=  "00000001111101";
		Trees_din <= x"040e6408";
		wait for Clk_period;
		Addr <=  "00000001111110";
		Trees_din <= x"06f48004";
		wait for Clk_period;
		Addr <=  "00000001111111";
		Trees_din <= x"ff840249";
		wait for Clk_period;
		Addr <=  "00000010000000";
		Trees_din <= x"009f0249";
		wait for Clk_period;
		Addr <=  "00000010000001";
		Trees_din <= x"017d0249";
		wait for Clk_period;
		Addr <=  "00000010000010";
		Trees_din <= x"1b003004";
		wait for Clk_period;
		Addr <=  "00000010000011";
		Trees_din <= x"01190249";
		wait for Clk_period;
		Addr <=  "00000010000100";
		Trees_din <= x"05f7cc04";
		wait for Clk_period;
		Addr <=  "00000010000101";
		Trees_din <= x"00930249";
		wait for Clk_period;
		Addr <=  "00000010000110";
		Trees_din <= x"ff600249";
		wait for Clk_period;
		Addr <=  "00000010000111";
		Trees_din <= x"19007f04";
		wait for Clk_period;
		Addr <=  "00000010001000";
		Trees_din <= x"01320249";
		wait for Clk_period;
		Addr <=  "00000010001001";
		Trees_din <= x"0e03c410";
		wait for Clk_period;
		Addr <=  "00000010001010";
		Trees_din <= x"10f95e08";
		wait for Clk_period;
		Addr <=  "00000010001011";
		Trees_din <= x"1b003b04";
		wait for Clk_period;
		Addr <=  "00000010001100";
		Trees_din <= x"ff990249";
		wait for Clk_period;
		Addr <=  "00000010001101";
		Trees_din <= x"00d70249";
		wait for Clk_period;
		Addr <=  "00000010001110";
		Trees_din <= x"15007f04";
		wait for Clk_period;
		Addr <=  "00000010001111";
		Trees_din <= x"00390249";
		wait for Clk_period;
		Addr <=  "00000010010000";
		Trees_din <= x"ff600249";
		wait for Clk_period;
		Addr <=  "00000010010001";
		Trees_din <= x"00b60249";
		wait for Clk_period;
		Addr <=  "00000010010010";
		Trees_din <= x"0406be5c";
		wait for Clk_period;
		Addr <=  "00000010010011";
		Trees_din <= x"04041b2c";
		wait for Clk_period;
		Addr <=  "00000010010100";
		Trees_din <= x"0401dd14";
		wait for Clk_period;
		Addr <=  "00000010010101";
		Trees_din <= x"03fbf604";
		wait for Clk_period;
		Addr <=  "00000010010110";
		Trees_din <= x"ff5903b5";
		wait for Clk_period;
		Addr <=  "00000010010111";
		Trees_din <= x"0e045b08";
		wait for Clk_period;
		Addr <=  "00000010011000";
		Trees_din <= x"0f03fb04";
		wait for Clk_period;
		Addr <=  "00000010011001";
		Trees_din <= x"ff5f03b5";
		wait for Clk_period;
		Addr <=  "00000010011010";
		Trees_din <= x"ffee03b5";
		wait for Clk_period;
		Addr <=  "00000010011011";
		Trees_din <= x"0bfb0104";
		wait for Clk_period;
		Addr <=  "00000010011100";
		Trees_din <= x"009e03b5";
		wait for Clk_period;
		Addr <=  "00000010011101";
		Trees_din <= x"ff7003b5";
		wait for Clk_period;
		Addr <=  "00000010011110";
		Trees_din <= x"06f5ff08";
		wait for Clk_period;
		Addr <=  "00000010011111";
		Trees_din <= x"15007c04";
		wait for Clk_period;
		Addr <=  "00000010100000";
		Trees_din <= x"003203b5";
		wait for Clk_period;
		Addr <=  "00000010100001";
		Trees_din <= x"ff5b03b5";
		wait for Clk_period;
		Addr <=  "00000010100010";
		Trees_din <= x"02041d08";
		wait for Clk_period;
		Addr <=  "00000010100011";
		Trees_din <= x"03041704";
		wait for Clk_period;
		Addr <=  "00000010100100";
		Trees_din <= x"ffe303b5";
		wait for Clk_period;
		Addr <=  "00000010100101";
		Trees_din <= x"ff6303b5";
		wait for Clk_period;
		Addr <=  "00000010100110";
		Trees_din <= x"09005404";
		wait for Clk_period;
		Addr <=  "00000010100111";
		Trees_din <= x"016603b5";
		wait for Clk_period;
		Addr <=  "00000010101000";
		Trees_din <= x"003903b5";
		wait for Clk_period;
		Addr <=  "00000010101001";
		Trees_din <= x"05fe311c";
		wait for Clk_period;
		Addr <=  "00000010101010";
		Trees_din <= x"0d03a510";
		wait for Clk_period;
		Addr <=  "00000010101011";
		Trees_din <= x"0c03a408";
		wait for Clk_period;
		Addr <=  "00000010101100";
		Trees_din <= x"1200f704";
		wait for Clk_period;
		Addr <=  "00000010101101";
		Trees_din <= x"ffeb03b5";
		wait for Clk_period;
		Addr <=  "00000010101110";
		Trees_din <= x"ff7603b5";
		wait for Clk_period;
		Addr <=  "00000010101111";
		Trees_din <= x"12032a04";
		wait for Clk_period;
		Addr <=  "00000010110000";
		Trees_din <= x"00b703b5";
		wait for Clk_period;
		Addr <=  "00000010110001";
		Trees_din <= x"ff9b03b5";
		wait for Clk_period;
		Addr <=  "00000010110010";
		Trees_din <= x"05faab04";
		wait for Clk_period;
		Addr <=  "00000010110011";
		Trees_din <= x"ff9003b5";
		wait for Clk_period;
		Addr <=  "00000010110100";
		Trees_din <= x"09005304";
		wait for Clk_period;
		Addr <=  "00000010110101";
		Trees_din <= x"017203b5";
		wait for Clk_period;
		Addr <=  "00000010110110";
		Trees_din <= x"001203b5";
		wait for Clk_period;
		Addr <=  "00000010110111";
		Trees_din <= x"0d02700c";
		wait for Clk_period;
		Addr <=  "00000010111000";
		Trees_din <= x"11026a04";
		wait for Clk_period;
		Addr <=  "00000010111001";
		Trees_din <= x"ff7d03b5";
		wait for Clk_period;
		Addr <=  "00000010111010";
		Trees_din <= x"11028704";
		wait for Clk_period;
		Addr <=  "00000010111011";
		Trees_din <= x"00fd03b5";
		wait for Clk_period;
		Addr <=  "00000010111100";
		Trees_din <= x"ff9b03b5";
		wait for Clk_period;
		Addr <=  "00000010111101";
		Trees_din <= x"0bf95804";
		wait for Clk_period;
		Addr <=  "00000010111110";
		Trees_din <= x"ff9b03b5";
		wait for Clk_period;
		Addr <=  "00000010111111";
		Trees_din <= x"017403b5";
		wait for Clk_period;
		Addr <=  "00000011000000";
		Trees_din <= x"040a4a34";
		wait for Clk_period;
		Addr <=  "00000011000001";
		Trees_din <= x"05fcf118";
		wait for Clk_period;
		Addr <=  "00000011000010";
		Trees_din <= x"09005910";
		wait for Clk_period;
		Addr <=  "00000011000011";
		Trees_din <= x"04077808";
		wait for Clk_period;
		Addr <=  "00000011000100";
		Trees_din <= x"1b003304";
		wait for Clk_period;
		Addr <=  "00000011000101";
		Trees_din <= x"007703b5";
		wait for Clk_period;
		Addr <=  "00000011000110";
		Trees_din <= x"ff5e03b5";
		wait for Clk_period;
		Addr <=  "00000011000111";
		Trees_din <= x"06f3ca04";
		wait for Clk_period;
		Addr <=  "00000011001000";
		Trees_din <= x"000003b5";
		wait for Clk_period;
		Addr <=  "00000011001001";
		Trees_din <= x"00c703b5";
		wait for Clk_period;
		Addr <=  "00000011001010";
		Trees_din <= x"0bf94a04";
		wait for Clk_period;
		Addr <=  "00000011001011";
		Trees_din <= x"00a603b5";
		wait for Clk_period;
		Addr <=  "00000011001100";
		Trees_din <= x"ff5903b5";
		wait for Clk_period;
		Addr <=  "00000011001101";
		Trees_din <= x"06f5850c";
		wait for Clk_period;
		Addr <=  "00000011001110";
		Trees_din <= x"0d023404";
		wait for Clk_period;
		Addr <=  "00000011001111";
		Trees_din <= x"ff6f03b5";
		wait for Clk_period;
		Addr <=  "00000011010000";
		Trees_din <= x"1401c004";
		wait for Clk_period;
		Addr <=  "00000011010001";
		Trees_din <= x"fff203b5";
		wait for Clk_period;
		Addr <=  "00000011010010";
		Trees_din <= x"010503b5";
		wait for Clk_period;
		Addr <=  "00000011010011";
		Trees_din <= x"1603ed08";
		wait for Clk_period;
		Addr <=  "00000011010100";
		Trees_din <= x"1d003904";
		wait for Clk_period;
		Addr <=  "00000011010101";
		Trees_din <= x"002303b5";
		wait for Clk_period;
		Addr <=  "00000011010110";
		Trees_din <= x"015603b5";
		wait for Clk_period;
		Addr <=  "00000011010111";
		Trees_din <= x"08004004";
		wait for Clk_period;
		Addr <=  "00000011011000";
		Trees_din <= x"009a03b5";
		wait for Clk_period;
		Addr <=  "00000011011001";
		Trees_din <= x"ff8b03b5";
		wait for Clk_period;
		Addr <=  "00000011011010";
		Trees_din <= x"03096514";
		wait for Clk_period;
		Addr <=  "00000011011011";
		Trees_din <= x"0ef8c504";
		wait for Clk_period;
		Addr <=  "00000011011100";
		Trees_din <= x"fff203b5";
		wait for Clk_period;
		Addr <=  "00000011011101";
		Trees_din <= x"02055108";
		wait for Clk_period;
		Addr <=  "00000011011110";
		Trees_din <= x"0e06a204";
		wait for Clk_period;
		Addr <=  "00000011011111";
		Trees_din <= x"013003b5";
		wait for Clk_period;
		Addr <=  "00000011100000";
		Trees_din <= x"fffe03b5";
		wait for Clk_period;
		Addr <=  "00000011100001";
		Trees_din <= x"01059504";
		wait for Clk_period;
		Addr <=  "00000011100010";
		Trees_din <= x"ff9c03b5";
		wait for Clk_period;
		Addr <=  "00000011100011";
		Trees_din <= x"00c803b5";
		wait for Clk_period;
		Addr <=  "00000011100100";
		Trees_din <= x"0f01080c";
		wait for Clk_period;
		Addr <=  "00000011100101";
		Trees_din <= x"10044d08";
		wait for Clk_period;
		Addr <=  "00000011100110";
		Trees_din <= x"0b026f04";
		wait for Clk_period;
		Addr <=  "00000011100111";
		Trees_din <= x"005903b5";
		wait for Clk_period;
		Addr <=  "00000011101000";
		Trees_din <= x"01bf03b5";
		wait for Clk_period;
		Addr <=  "00000011101001";
		Trees_din <= x"ffe903b5";
		wait for Clk_period;
		Addr <=  "00000011101010";
		Trees_din <= x"02001704";
		wait for Clk_period;
		Addr <=  "00000011101011";
		Trees_din <= x"ff6903b5";
		wait for Clk_period;
		Addr <=  "00000011101100";
		Trees_din <= x"002303b5";
		wait for Clk_period;
		Addr <=  "00000011101101";
		Trees_din <= x"04045e48";
		wait for Clk_period;
		Addr <=  "00000011101110";
		Trees_din <= x"0401dd20";
		wait for Clk_period;
		Addr <=  "00000011101111";
		Trees_din <= x"03fbf604";
		wait for Clk_period;
		Addr <=  "00000011110000";
		Trees_din <= x"ff5c04d9";
		wait for Clk_period;
		Addr <=  "00000011110001";
		Trees_din <= x"0e045b10";
		wait for Clk_period;
		Addr <=  "00000011110010";
		Trees_din <= x"0c004308";
		wait for Clk_period;
		Addr <=  "00000011110011";
		Trees_din <= x"1b003604";
		wait for Clk_period;
		Addr <=  "00000011110100";
		Trees_din <= x"011504d9";
		wait for Clk_period;
		Addr <=  "00000011110101";
		Trees_din <= x"ff6f04d9";
		wait for Clk_period;
		Addr <=  "00000011110110";
		Trees_din <= x"09003c04";
		wait for Clk_period;
		Addr <=  "00000011110111";
		Trees_din <= x"002404d9";
		wait for Clk_period;
		Addr <=  "00000011111000";
		Trees_din <= x"ff6004d9";
		wait for Clk_period;
		Addr <=  "00000011111001";
		Trees_din <= x"0bfb0108";
		wait for Clk_period;
		Addr <=  "00000011111010";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00000011111011";
		Trees_din <= x"017004d9";
		wait for Clk_period;
		Addr <=  "00000011111100";
		Trees_din <= x"ff9b04d9";
		wait for Clk_period;
		Addr <=  "00000011111101";
		Trees_din <= x"ff7804d9";
		wait for Clk_period;
		Addr <=  "00000011111110";
		Trees_din <= x"0efcb010";
		wait for Clk_period;
		Addr <=  "00000011111111";
		Trees_din <= x"16009a04";
		wait for Clk_period;
		Addr <=  "00000100000000";
		Trees_din <= x"ff7c04d9";
		wait for Clk_period;
		Addr <=  "00000100000001";
		Trees_din <= x"00ff2d04";
		wait for Clk_period;
		Addr <=  "00000100000010";
		Trees_din <= x"ff9904d9";
		wait for Clk_period;
		Addr <=  "00000100000011";
		Trees_din <= x"1a00cc04";
		wait for Clk_period;
		Addr <=  "00000100000100";
		Trees_din <= x"019304d9";
		wait for Clk_period;
		Addr <=  "00000100000101";
		Trees_din <= x"002f04d9";
		wait for Clk_period;
		Addr <=  "00000100000110";
		Trees_din <= x"04025d0c";
		wait for Clk_period;
		Addr <=  "00000100000111";
		Trees_din <= x"06f5ff04";
		wait for Clk_period;
		Addr <=  "00000100001000";
		Trees_din <= x"ff7604d9";
		wait for Clk_period;
		Addr <=  "00000100001001";
		Trees_din <= x"02ffb904";
		wait for Clk_period;
		Addr <=  "00000100001010";
		Trees_din <= x"ff8504d9";
		wait for Clk_period;
		Addr <=  "00000100001011";
		Trees_din <= x"014504d9";
		wait for Clk_period;
		Addr <=  "00000100001100";
		Trees_din <= x"05feb404";
		wait for Clk_period;
		Addr <=  "00000100001101";
		Trees_din <= x"ff5d04d9";
		wait for Clk_period;
		Addr <=  "00000100001110";
		Trees_din <= x"11029c04";
		wait for Clk_period;
		Addr <=  "00000100001111";
		Trees_din <= x"ff8204d9";
		wait for Clk_period;
		Addr <=  "00000100010000";
		Trees_din <= x"003904d9";
		wait for Clk_period;
		Addr <=  "00000100010001";
		Trees_din <= x"0409d634";
		wait for Clk_period;
		Addr <=  "00000100010010";
		Trees_din <= x"05fcd01c";
		wait for Clk_period;
		Addr <=  "00000100010011";
		Trees_din <= x"0d03a50c";
		wait for Clk_period;
		Addr <=  "00000100010100";
		Trees_din <= x"1104d508";
		wait for Clk_period;
		Addr <=  "00000100010101";
		Trees_din <= x"16000504";
		wait for Clk_period;
		Addr <=  "00000100010110";
		Trees_din <= x"009d04d9";
		wait for Clk_period;
		Addr <=  "00000100010111";
		Trees_din <= x"ffc304d9";
		wait for Clk_period;
		Addr <=  "00000100011000";
		Trees_din <= x"012c04d9";
		wait for Clk_period;
		Addr <=  "00000100011001";
		Trees_din <= x"06f56508";
		wait for Clk_period;
		Addr <=  "00000100011010";
		Trees_din <= x"06f2a604";
		wait for Clk_period;
		Addr <=  "00000100011011";
		Trees_din <= x"000f04d9";
		wait for Clk_period;
		Addr <=  "00000100011100";
		Trees_din <= x"019604d9";
		wait for Clk_period;
		Addr <=  "00000100011101";
		Trees_din <= x"07005a04";
		wait for Clk_period;
		Addr <=  "00000100011110";
		Trees_din <= x"003304d9";
		wait for Clk_period;
		Addr <=  "00000100011111";
		Trees_din <= x"ff9704d9";
		wait for Clk_period;
		Addr <=  "00000100100000";
		Trees_din <= x"06f5720c";
		wait for Clk_period;
		Addr <=  "00000100100001";
		Trees_din <= x"0d023404";
		wait for Clk_period;
		Addr <=  "00000100100010";
		Trees_din <= x"ff6904d9";
		wait for Clk_period;
		Addr <=  "00000100100011";
		Trees_din <= x"0204f604";
		wait for Clk_period;
		Addr <=  "00000100100100";
		Trees_din <= x"00b604d9";
		wait for Clk_period;
		Addr <=  "00000100100101";
		Trees_din <= x"ff8704d9";
		wait for Clk_period;
		Addr <=  "00000100100110";
		Trees_din <= x"1d003804";
		wait for Clk_period;
		Addr <=  "00000100100111";
		Trees_din <= x"ff7204d9";
		wait for Clk_period;
		Addr <=  "00000100101000";
		Trees_din <= x"14004f04";
		wait for Clk_period;
		Addr <=  "00000100101001";
		Trees_din <= x"ffcf04d9";
		wait for Clk_period;
		Addr <=  "00000100101010";
		Trees_din <= x"00d204d9";
		wait for Clk_period;
		Addr <=  "00000100101011";
		Trees_din <= x"040e6414";
		wait for Clk_period;
		Addr <=  "00000100101100";
		Trees_din <= x"05f7b504";
		wait for Clk_period;
		Addr <=  "00000100101101";
		Trees_din <= x"ff7304d9";
		wait for Clk_period;
		Addr <=  "00000100101110";
		Trees_din <= x"01074708";
		wait for Clk_period;
		Addr <=  "00000100101111";
		Trees_din <= x"1005b204";
		wait for Clk_period;
		Addr <=  "00000100110000";
		Trees_din <= x"00cd04d9";
		wait for Clk_period;
		Addr <=  "00000100110001";
		Trees_din <= x"ffae04d9";
		wait for Clk_period;
		Addr <=  "00000100110010";
		Trees_din <= x"12029604";
		wait for Clk_period;
		Addr <=  "00000100110011";
		Trees_din <= x"ff8a04d9";
		wait for Clk_period;
		Addr <=  "00000100110100";
		Trees_din <= x"00fd04d9";
		wait for Clk_period;
		Addr <=  "00000100110101";
		Trees_din <= x"011204d9";
		wait for Clk_period;
		Addr <=  "00000100110110";
		Trees_din <= x"04045e3c";
		wait for Clk_period;
		Addr <=  "00000100110111";
		Trees_din <= x"04007b18";
		wait for Clk_period;
		Addr <=  "00000100111000";
		Trees_din <= x"0e045b0c";
		wait for Clk_period;
		Addr <=  "00000100111001";
		Trees_din <= x"0215a804";
		wait for Clk_period;
		Addr <=  "00000100111010";
		Trees_din <= x"ff5f05dd";
		wait for Clk_period;
		Addr <=  "00000100111011";
		Trees_din <= x"1a00a304";
		wait for Clk_period;
		Addr <=  "00000100111100";
		Trees_din <= x"004805dd";
		wait for Clk_period;
		Addr <=  "00000100111101";
		Trees_din <= x"ff7a05dd";
		wait for Clk_period;
		Addr <=  "00000100111110";
		Trees_din <= x"03fce704";
		wait for Clk_period;
		Addr <=  "00000100111111";
		Trees_din <= x"ff6405dd";
		wait for Clk_period;
		Addr <=  "00000101000000";
		Trees_din <= x"11043104";
		wait for Clk_period;
		Addr <=  "00000101000001";
		Trees_din <= x"ff8805dd";
		wait for Clk_period;
		Addr <=  "00000101000010";
		Trees_din <= x"00eb05dd";
		wait for Clk_period;
		Addr <=  "00000101000011";
		Trees_din <= x"10052d10";
		wait for Clk_period;
		Addr <=  "00000101000100";
		Trees_din <= x"0d000004";
		wait for Clk_period;
		Addr <=  "00000101000101";
		Trees_din <= x"006b05dd";
		wait for Clk_period;
		Addr <=  "00000101000110";
		Trees_din <= x"0a077008";
		wait for Clk_period;
		Addr <=  "00000101000111";
		Trees_din <= x"0ef99404";
		wait for Clk_period;
		Addr <=  "00000101001000";
		Trees_din <= x"ffce05dd";
		wait for Clk_period;
		Addr <=  "00000101001001";
		Trees_din <= x"ff6905dd";
		wait for Clk_period;
		Addr <=  "00000101001010";
		Trees_din <= x"003a05dd";
		wait for Clk_period;
		Addr <=  "00000101001011";
		Trees_din <= x"19009e08";
		wait for Clk_period;
		Addr <=  "00000101001100";
		Trees_din <= x"05f8b404";
		wait for Clk_period;
		Addr <=  "00000101001101";
		Trees_din <= x"003d05dd";
		wait for Clk_period;
		Addr <=  "00000101001110";
		Trees_din <= x"ff6e05dd";
		wait for Clk_period;
		Addr <=  "00000101001111";
		Trees_din <= x"0c01d304";
		wait for Clk_period;
		Addr <=  "00000101010000";
		Trees_din <= x"ff8d05dd";
		wait for Clk_period;
		Addr <=  "00000101010001";
		Trees_din <= x"1200ae04";
		wait for Clk_period;
		Addr <=  "00000101010010";
		Trees_din <= x"001f05dd";
		wait for Clk_period;
		Addr <=  "00000101010011";
		Trees_din <= x"016405dd";
		wait for Clk_period;
		Addr <=  "00000101010100";
		Trees_din <= x"0409d624";
		wait for Clk_period;
		Addr <=  "00000101010101";
		Trees_din <= x"07004d04";
		wait for Clk_period;
		Addr <=  "00000101010110";
		Trees_din <= x"ff6605dd";
		wait for Clk_period;
		Addr <=  "00000101010111";
		Trees_din <= x"09005310";
		wait for Clk_period;
		Addr <=  "00000101011000";
		Trees_din <= x"0d039d08";
		wait for Clk_period;
		Addr <=  "00000101011001";
		Trees_din <= x"05fb5604";
		wait for Clk_period;
		Addr <=  "00000101011010";
		Trees_din <= x"ffbb05dd";
		wait for Clk_period;
		Addr <=  "00000101011011";
		Trees_din <= x"008105dd";
		wait for Clk_period;
		Addr <=  "00000101011100";
		Trees_din <= x"01fdac04";
		wait for Clk_period;
		Addr <=  "00000101011101";
		Trees_din <= x"005105dd";
		wait for Clk_period;
		Addr <=  "00000101011110";
		Trees_din <= x"015605dd";
		wait for Clk_period;
		Addr <=  "00000101011111";
		Trees_din <= x"17000008";
		wait for Clk_period;
		Addr <=  "00000101100000";
		Trees_din <= x"0406be04";
		wait for Clk_period;
		Addr <=  "00000101100001";
		Trees_din <= x"ffec05dd";
		wait for Clk_period;
		Addr <=  "00000101100010";
		Trees_din <= x"00a005dd";
		wait for Clk_period;
		Addr <=  "00000101100011";
		Trees_din <= x"05fcf104";
		wait for Clk_period;
		Addr <=  "00000101100100";
		Trees_din <= x"ff9505dd";
		wait for Clk_period;
		Addr <=  "00000101100101";
		Trees_din <= x"001f05dd";
		wait for Clk_period;
		Addr <=  "00000101100110";
		Trees_din <= x"040e6414";
		wait for Clk_period;
		Addr <=  "00000101100111";
		Trees_din <= x"05f7b504";
		wait for Clk_period;
		Addr <=  "00000101101000";
		Trees_din <= x"ff7b05dd";
		wait for Clk_period;
		Addr <=  "00000101101001";
		Trees_din <= x"0bf9ce08";
		wait for Clk_period;
		Addr <=  "00000101101010";
		Trees_din <= x"11029704";
		wait for Clk_period;
		Addr <=  "00000101101011";
		Trees_din <= x"ff5605dd";
		wait for Clk_period;
		Addr <=  "00000101101100";
		Trees_din <= x"008205dd";
		wait for Clk_period;
		Addr <=  "00000101101101";
		Trees_din <= x"07005e04";
		wait for Clk_period;
		Addr <=  "00000101101110";
		Trees_din <= x"00a405dd";
		wait for Clk_period;
		Addr <=  "00000101101111";
		Trees_din <= x"ff7305dd";
		wait for Clk_period;
		Addr <=  "00000101110000";
		Trees_din <= x"12fbf704";
		wait for Clk_period;
		Addr <=  "00000101110001";
		Trees_din <= x"000b05dd";
		wait for Clk_period;
		Addr <=  "00000101110010";
		Trees_din <= x"0bf96508";
		wait for Clk_period;
		Addr <=  "00000101110011";
		Trees_din <= x"09005504";
		wait for Clk_period;
		Addr <=  "00000101110100";
		Trees_din <= x"ffcf05dd";
		wait for Clk_period;
		Addr <=  "00000101110101";
		Trees_din <= x"00d005dd";
		wait for Clk_period;
		Addr <=  "00000101110110";
		Trees_din <= x"00fd05dd";
		wait for Clk_period;
		Addr <=  "00000101110111";
		Trees_din <= x"04045e48";
		wait for Clk_period;
		Addr <=  "00000101111000";
		Trees_din <= x"04007b20";
		wait for Clk_period;
		Addr <=  "00000101111001";
		Trees_din <= x"0e045b14";
		wait for Clk_period;
		Addr <=  "00000101111010";
		Trees_din <= x"0215a80c";
		wait for Clk_period;
		Addr <=  "00000101111011";
		Trees_din <= x"09003c08";
		wait for Clk_period;
		Addr <=  "00000101111100";
		Trees_din <= x"08015304";
		wait for Clk_period;
		Addr <=  "00000101111101";
		Trees_din <= x"ff7906d9";
		wait for Clk_period;
		Addr <=  "00000101111110";
		Trees_din <= x"004506d9";
		wait for Clk_period;
		Addr <=  "00000101111111";
		Trees_din <= x"ff6106d9";
		wait for Clk_period;
		Addr <=  "00000110000000";
		Trees_din <= x"1e007604";
		wait for Clk_period;
		Addr <=  "00000110000001";
		Trees_din <= x"ff8106d9";
		wait for Clk_period;
		Addr <=  "00000110000010";
		Trees_din <= x"004406d9";
		wait for Clk_period;
		Addr <=  "00000110000011";
		Trees_din <= x"03fce704";
		wait for Clk_period;
		Addr <=  "00000110000100";
		Trees_din <= x"ff6706d9";
		wait for Clk_period;
		Addr <=  "00000110000101";
		Trees_din <= x"11043104";
		wait for Clk_period;
		Addr <=  "00000110000110";
		Trees_din <= x"ff8f06d9";
		wait for Clk_period;
		Addr <=  "00000110000111";
		Trees_din <= x"00c906d9";
		wait for Clk_period;
		Addr <=  "00000110001000";
		Trees_din <= x"05fe7018";
		wait for Clk_period;
		Addr <=  "00000110001001";
		Trees_din <= x"0d000408";
		wait for Clk_period;
		Addr <=  "00000110001010";
		Trees_din <= x"0c004104";
		wait for Clk_period;
		Addr <=  "00000110001011";
		Trees_din <= x"00ce06d9";
		wait for Clk_period;
		Addr <=  "00000110001100";
		Trees_din <= x"ff8906d9";
		wait for Clk_period;
		Addr <=  "00000110001101";
		Trees_din <= x"0f000c08";
		wait for Clk_period;
		Addr <=  "00000110001110";
		Trees_din <= x"14012a04";
		wait for Clk_period;
		Addr <=  "00000110001111";
		Trees_din <= x"ff7906d9";
		wait for Clk_period;
		Addr <=  "00000110010000";
		Trees_din <= x"009e06d9";
		wait for Clk_period;
		Addr <=  "00000110010001";
		Trees_din <= x"1a008d04";
		wait for Clk_period;
		Addr <=  "00000110010010";
		Trees_din <= x"001d06d9";
		wait for Clk_period;
		Addr <=  "00000110010011";
		Trees_din <= x"ff6806d9";
		wait for Clk_period;
		Addr <=  "00000110010100";
		Trees_din <= x"10052508";
		wait for Clk_period;
		Addr <=  "00000110010101";
		Trees_din <= x"0efb0d04";
		wait for Clk_period;
		Addr <=  "00000110010110";
		Trees_din <= x"005506d9";
		wait for Clk_period;
		Addr <=  "00000110010111";
		Trees_din <= x"ff7006d9";
		wait for Clk_period;
		Addr <=  "00000110011000";
		Trees_din <= x"19009d04";
		wait for Clk_period;
		Addr <=  "00000110011001";
		Trees_din <= x"ff9d06d9";
		wait for Clk_period;
		Addr <=  "00000110011010";
		Trees_din <= x"011306d9";
		wait for Clk_period;
		Addr <=  "00000110011011";
		Trees_din <= x"040e6428";
		wait for Clk_period;
		Addr <=  "00000110011100";
		Trees_din <= x"07005614";
		wait for Clk_period;
		Addr <=  "00000110011101";
		Trees_din <= x"06f1ee04";
		wait for Clk_period;
		Addr <=  "00000110011110";
		Trees_din <= x"ff7406d9";
		wait for Clk_period;
		Addr <=  "00000110011111";
		Trees_din <= x"1900a908";
		wait for Clk_period;
		Addr <=  "00000110100000";
		Trees_din <= x"19009b04";
		wait for Clk_period;
		Addr <=  "00000110100001";
		Trees_din <= x"005806d9";
		wait for Clk_period;
		Addr <=  "00000110100010";
		Trees_din <= x"00d306d9";
		wait for Clk_period;
		Addr <=  "00000110100011";
		Trees_din <= x"0afe5a04";
		wait for Clk_period;
		Addr <=  "00000110100100";
		Trees_din <= x"ffbd06d9";
		wait for Clk_period;
		Addr <=  "00000110100101";
		Trees_din <= x"005d06d9";
		wait for Clk_period;
		Addr <=  "00000110100110";
		Trees_din <= x"1104d510";
		wait for Clk_period;
		Addr <=  "00000110100111";
		Trees_din <= x"06f45808";
		wait for Clk_period;
		Addr <=  "00000110101000";
		Trees_din <= x"0af7ba04";
		wait for Clk_period;
		Addr <=  "00000110101001";
		Trees_din <= x"00af06d9";
		wait for Clk_period;
		Addr <=  "00000110101010";
		Trees_din <= x"ffaa06d9";
		wait for Clk_period;
		Addr <=  "00000110101011";
		Trees_din <= x"1500a004";
		wait for Clk_period;
		Addr <=  "00000110101100";
		Trees_din <= x"000e06d9";
		wait for Clk_period;
		Addr <=  "00000110101101";
		Trees_din <= x"009406d9";
		wait for Clk_period;
		Addr <=  "00000110101110";
		Trees_din <= x"011f06d9";
		wait for Clk_period;
		Addr <=  "00000110101111";
		Trees_din <= x"12fbf704";
		wait for Clk_period;
		Addr <=  "00000110110000";
		Trees_din <= x"000806d9";
		wait for Clk_period;
		Addr <=  "00000110110001";
		Trees_din <= x"0bf96508";
		wait for Clk_period;
		Addr <=  "00000110110010";
		Trees_din <= x"09005504";
		wait for Clk_period;
		Addr <=  "00000110110011";
		Trees_din <= x"ffd106d9";
		wait for Clk_period;
		Addr <=  "00000110110100";
		Trees_din <= x"00ba06d9";
		wait for Clk_period;
		Addr <=  "00000110110101";
		Trees_din <= x"00df06d9";
		wait for Clk_period;
		Addr <=  "00000110110110";
		Trees_din <= x"04045e3c";
		wait for Clk_period;
		Addr <=  "00000110110111";
		Trees_din <= x"04007b20";
		wait for Clk_period;
		Addr <=  "00000110111000";
		Trees_din <= x"0e045b14";
		wait for Clk_period;
		Addr <=  "00000110111001";
		Trees_din <= x"0215a80c";
		wait for Clk_period;
		Addr <=  "00000110111010";
		Trees_din <= x"09003c08";
		wait for Clk_period;
		Addr <=  "00000110111011";
		Trees_din <= x"17000004";
		wait for Clk_period;
		Addr <=  "00000110111100";
		Trees_din <= x"004807f5";
		wait for Clk_period;
		Addr <=  "00000110111101";
		Trees_din <= x"ff7f07f5";
		wait for Clk_period;
		Addr <=  "00000110111110";
		Trees_din <= x"ff6307f5";
		wait for Clk_period;
		Addr <=  "00000110111111";
		Trees_din <= x"1603e504";
		wait for Clk_period;
		Addr <=  "00000111000000";
		Trees_din <= x"ff8807f5";
		wait for Clk_period;
		Addr <=  "00000111000001";
		Trees_din <= x"004907f5";
		wait for Clk_period;
		Addr <=  "00000111000010";
		Trees_din <= x"03fce704";
		wait for Clk_period;
		Addr <=  "00000111000011";
		Trees_din <= x"ff6a07f5";
		wait for Clk_period;
		Addr <=  "00000111000100";
		Trees_din <= x"0bfb0104";
		wait for Clk_period;
		Addr <=  "00000111000101";
		Trees_din <= x"00bb07f5";
		wait for Clk_period;
		Addr <=  "00000111000110";
		Trees_din <= x"ff9407f5";
		wait for Clk_period;
		Addr <=  "00000111000111";
		Trees_din <= x"06f4ea04";
		wait for Clk_period;
		Addr <=  "00000111001000";
		Trees_din <= x"ff6707f5";
		wait for Clk_period;
		Addr <=  "00000111001001";
		Trees_din <= x"02ff8608";
		wait for Clk_period;
		Addr <=  "00000111001010";
		Trees_din <= x"0b053004";
		wait for Clk_period;
		Addr <=  "00000111001011";
		Trees_din <= x"ff6a07f5";
		wait for Clk_period;
		Addr <=  "00000111001100";
		Trees_din <= x"fff307f5";
		wait for Clk_period;
		Addr <=  "00000111001101";
		Trees_din <= x"0b036f08";
		wait for Clk_period;
		Addr <=  "00000111001110";
		Trees_din <= x"1a00be04";
		wait for Clk_period;
		Addr <=  "00000111001111";
		Trees_din <= x"ffcf07f5";
		wait for Clk_period;
		Addr <=  "00000111010000";
		Trees_din <= x"00a107f5";
		wait for Clk_period;
		Addr <=  "00000111010001";
		Trees_din <= x"10f74f04";
		wait for Clk_period;
		Addr <=  "00000111010010";
		Trees_din <= x"002e07f5";
		wait for Clk_period;
		Addr <=  "00000111010011";
		Trees_din <= x"ff7007f5";
		wait for Clk_period;
		Addr <=  "00000111010100";
		Trees_din <= x"0409d624";
		wait for Clk_period;
		Addr <=  "00000111010101";
		Trees_din <= x"07004d04";
		wait for Clk_period;
		Addr <=  "00000111010110";
		Trees_din <= x"ff6a07f5";
		wait for Clk_period;
		Addr <=  "00000111010111";
		Trees_din <= x"09005310";
		wait for Clk_period;
		Addr <=  "00000111011000";
		Trees_din <= x"0d039d08";
		wait for Clk_period;
		Addr <=  "00000111011001";
		Trees_din <= x"0308a904";
		wait for Clk_period;
		Addr <=  "00000111011010";
		Trees_din <= x"005007f5";
		wait for Clk_period;
		Addr <=  "00000111011011";
		Trees_din <= x"ff9807f5";
		wait for Clk_period;
		Addr <=  "00000111011100";
		Trees_din <= x"1a00b604";
		wait for Clk_period;
		Addr <=  "00000111011101";
		Trees_din <= x"005f07f5";
		wait for Clk_period;
		Addr <=  "00000111011110";
		Trees_din <= x"012907f5";
		wait for Clk_period;
		Addr <=  "00000111011111";
		Trees_din <= x"1400eb08";
		wait for Clk_period;
		Addr <=  "00000111100000";
		Trees_din <= x"0c003204";
		wait for Clk_period;
		Addr <=  "00000111100001";
		Trees_din <= x"002207f5";
		wait for Clk_period;
		Addr <=  "00000111100010";
		Trees_din <= x"ff7407f5";
		wait for Clk_period;
		Addr <=  "00000111100011";
		Trees_din <= x"1104d504";
		wait for Clk_period;
		Addr <=  "00000111100100";
		Trees_din <= x"001807f5";
		wait for Clk_period;
		Addr <=  "00000111100101";
		Trees_din <= x"012107f5";
		wait for Clk_period;
		Addr <=  "00000111100110";
		Trees_din <= x"040e6420";
		wait for Clk_period;
		Addr <=  "00000111100111";
		Trees_din <= x"1a00d910";
		wait for Clk_period;
		Addr <=  "00000111101000";
		Trees_din <= x"0105dd08";
		wait for Clk_period;
		Addr <=  "00000111101001";
		Trees_din <= x"02023e04";
		wait for Clk_period;
		Addr <=  "00000111101010";
		Trees_din <= x"006f07f5";
		wait for Clk_period;
		Addr <=  "00000111101011";
		Trees_din <= x"ffa607f5";
		wait for Clk_period;
		Addr <=  "00000111101100";
		Trees_din <= x"11000d04";
		wait for Clk_period;
		Addr <=  "00000111101101";
		Trees_din <= x"003207f5";
		wait for Clk_period;
		Addr <=  "00000111101110";
		Trees_din <= x"ff5507f5";
		wait for Clk_period;
		Addr <=  "00000111101111";
		Trees_din <= x"03096508";
		wait for Clk_period;
		Addr <=  "00000111110000";
		Trees_din <= x"1703b604";
		wait for Clk_period;
		Addr <=  "00000111110001";
		Trees_din <= x"00c807f5";
		wait for Clk_period;
		Addr <=  "00000111110010";
		Trees_din <= x"ffb807f5";
		wait for Clk_period;
		Addr <=  "00000111110011";
		Trees_din <= x"1a00f904";
		wait for Clk_period;
		Addr <=  "00000111110100";
		Trees_din <= x"000c07f5";
		wait for Clk_period;
		Addr <=  "00000111110101";
		Trees_din <= x"ff8207f5";
		wait for Clk_period;
		Addr <=  "00000111110110";
		Trees_din <= x"12fbf704";
		wait for Clk_period;
		Addr <=  "00000111110111";
		Trees_din <= x"000707f5";
		wait for Clk_period;
		Addr <=  "00000111111000";
		Trees_din <= x"0bf96508";
		wait for Clk_period;
		Addr <=  "00000111111001";
		Trees_din <= x"09005504";
		wait for Clk_period;
		Addr <=  "00000111111010";
		Trees_din <= x"ffcf07f5";
		wait for Clk_period;
		Addr <=  "00000111111011";
		Trees_din <= x"00a607f5";
		wait for Clk_period;
		Addr <=  "00000111111100";
		Trees_din <= x"00ca07f5";
		wait for Clk_period;
		Addr <=  "00000111111101";
		Trees_din <= x"04041b40";
		wait for Clk_period;
		Addr <=  "00000111111110";
		Trees_din <= x"04fff320";
		wait for Clk_period;
		Addr <=  "00000111111111";
		Trees_din <= x"0215a818";
		wait for Clk_period;
		Addr <=  "00001000000000";
		Trees_din <= x"0e04b110";
		wait for Clk_period;
		Addr <=  "00001000000001";
		Trees_din <= x"09003c08";
		wait for Clk_period;
		Addr <=  "00001000000010";
		Trees_din <= x"0d039004";
		wait for Clk_period;
		Addr <=  "00001000000011";
		Trees_din <= x"ff860909";
		wait for Clk_period;
		Addr <=  "00001000000100";
		Trees_din <= x"00470909";
		wait for Clk_period;
		Addr <=  "00001000000101";
		Trees_din <= x"1703f604";
		wait for Clk_period;
		Addr <=  "00001000000110";
		Trees_din <= x"ff640909";
		wait for Clk_period;
		Addr <=  "00001000000111";
		Trees_din <= x"ffa20909";
		wait for Clk_period;
		Addr <=  "00001000001000";
		Trees_din <= x"04fd3f04";
		wait for Clk_period;
		Addr <=  "00001000001001";
		Trees_din <= x"ff720909";
		wait for Clk_period;
		Addr <=  "00001000001010";
		Trees_din <= x"005c0909";
		wait for Clk_period;
		Addr <=  "00001000001011";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00001000001100";
		Trees_din <= x"00480909";
		wait for Clk_period;
		Addr <=  "00001000001101";
		Trees_din <= x"ff8f0909";
		wait for Clk_period;
		Addr <=  "00001000001110";
		Trees_din <= x"06f5ff08";
		wait for Clk_period;
		Addr <=  "00001000001111";
		Trees_din <= x"18005104";
		wait for Clk_period;
		Addr <=  "00001000010000";
		Trees_din <= x"ff660909";
		wait for Clk_period;
		Addr <=  "00001000010001";
		Trees_din <= x"002f0909";
		wait for Clk_period;
		Addr <=  "00001000010010";
		Trees_din <= x"02ff7d08";
		wait for Clk_period;
		Addr <=  "00001000010011";
		Trees_din <= x"0b053004";
		wait for Clk_period;
		Addr <=  "00001000010100";
		Trees_din <= x"ff6e0909";
		wait for Clk_period;
		Addr <=  "00001000010101";
		Trees_din <= x"00030909";
		wait for Clk_period;
		Addr <=  "00001000010110";
		Trees_din <= x"0b028608";
		wait for Clk_period;
		Addr <=  "00001000010111";
		Trees_din <= x"1a00b804";
		wait for Clk_period;
		Addr <=  "00001000011000";
		Trees_din <= x"ff9c0909";
		wait for Clk_period;
		Addr <=  "00001000011001";
		Trees_din <= x"00b80909";
		wait for Clk_period;
		Addr <=  "00001000011010";
		Trees_din <= x"0f000f04";
		wait for Clk_period;
		Addr <=  "00001000011011";
		Trees_din <= x"00400909";
		wait for Clk_period;
		Addr <=  "00001000011100";
		Trees_din <= x"ff7d0909";
		wait for Clk_period;
		Addr <=  "00001000011101";
		Trees_din <= x"040e643c";
		wait for Clk_period;
		Addr <=  "00001000011110";
		Trees_din <= x"0406be1c";
		wait for Clk_period;
		Addr <=  "00001000011111";
		Trees_din <= x"11045610";
		wait for Clk_period;
		Addr <=  "00001000100000";
		Trees_din <= x"0f003708";
		wait for Clk_period;
		Addr <=  "00001000100001";
		Trees_din <= x"15009f04";
		wait for Clk_period;
		Addr <=  "00001000100010";
		Trees_din <= x"ffc60909";
		wait for Clk_period;
		Addr <=  "00001000100011";
		Trees_din <= x"00ca0909";
		wait for Clk_period;
		Addr <=  "00001000100100";
		Trees_din <= x"16000504";
		wait for Clk_period;
		Addr <=  "00001000100101";
		Trees_din <= x"007b0909";
		wait for Clk_period;
		Addr <=  "00001000100110";
		Trees_din <= x"ffa10909";
		wait for Clk_period;
		Addr <=  "00001000100111";
		Trees_din <= x"00fe7b04";
		wait for Clk_period;
		Addr <=  "00001000101000";
		Trees_din <= x"ffe10909";
		wait for Clk_period;
		Addr <=  "00001000101001";
		Trees_din <= x"08005c04";
		wait for Clk_period;
		Addr <=  "00001000101010";
		Trees_din <= x"01070909";
		wait for Clk_period;
		Addr <=  "00001000101011";
		Trees_din <= x"004e0909";
		wait for Clk_period;
		Addr <=  "00001000101100";
		Trees_din <= x"07005810";
		wait for Clk_period;
		Addr <=  "00001000101101";
		Trees_din <= x"01fd9408";
		wait for Clk_period;
		Addr <=  "00001000101110";
		Trees_din <= x"05fd7104";
		wait for Clk_period;
		Addr <=  "00001000101111";
		Trees_din <= x"00360909";
		wait for Clk_period;
		Addr <=  "00001000110000";
		Trees_din <= x"ff770909";
		wait for Clk_period;
		Addr <=  "00001000110001";
		Trees_din <= x"1a009f04";
		wait for Clk_period;
		Addr <=  "00001000110010";
		Trees_din <= x"ff7e0909";
		wait for Clk_period;
		Addr <=  "00001000110011";
		Trees_din <= x"007c0909";
		wait for Clk_period;
		Addr <=  "00001000110100";
		Trees_din <= x"11012208";
		wait for Clk_period;
		Addr <=  "00001000110101";
		Trees_din <= x"1e007404";
		wait for Clk_period;
		Addr <=  "00001000110110";
		Trees_din <= x"00000909";
		wait for Clk_period;
		Addr <=  "00001000110111";
		Trees_din <= x"00ed0909";
		wait for Clk_period;
		Addr <=  "00001000111000";
		Trees_din <= x"18004204";
		wait for Clk_period;
		Addr <=  "00001000111001";
		Trees_din <= x"002d0909";
		wait for Clk_period;
		Addr <=  "00001000111010";
		Trees_din <= x"ff9a0909";
		wait for Clk_period;
		Addr <=  "00001000111011";
		Trees_din <= x"12fbf704";
		wait for Clk_period;
		Addr <=  "00001000111100";
		Trees_din <= x"00080909";
		wait for Clk_period;
		Addr <=  "00001000111101";
		Trees_din <= x"0bf96508";
		wait for Clk_period;
		Addr <=  "00001000111110";
		Trees_din <= x"09005504";
		wait for Clk_period;
		Addr <=  "00001000111111";
		Trees_din <= x"ffd10909";
		wait for Clk_period;
		Addr <=  "00001001000000";
		Trees_din <= x"00990909";
		wait for Clk_period;
		Addr <=  "00001001000001";
		Trees_din <= x"00bb0909";
		wait for Clk_period;
		Addr <=  "00001001000010";
		Trees_din <= x"04041b34";
		wait for Clk_period;
		Addr <=  "00001001000011";
		Trees_din <= x"04fd5314";
		wait for Clk_period;
		Addr <=  "00001001000100";
		Trees_din <= x"0215a80c";
		wait for Clk_period;
		Addr <=  "00001001000101";
		Trees_din <= x"09003c08";
		wait for Clk_period;
		Addr <=  "00001001000110";
		Trees_din <= x"13fd7f04";
		wait for Clk_period;
		Addr <=  "00001001000111";
		Trees_din <= x"004509e5";
		wait for Clk_period;
		Addr <=  "00001001001000";
		Trees_din <= x"ff9309e5";
		wait for Clk_period;
		Addr <=  "00001001001001";
		Trees_din <= x"ff6409e5";
		wait for Clk_period;
		Addr <=  "00001001001010";
		Trees_din <= x"04fa8004";
		wait for Clk_period;
		Addr <=  "00001001001011";
		Trees_din <= x"ff9e09e5";
		wait for Clk_period;
		Addr <=  "00001001001100";
		Trees_din <= x"004709e5";
		wait for Clk_period;
		Addr <=  "00001001001101";
		Trees_din <= x"06f5ff08";
		wait for Clk_period;
		Addr <=  "00001001001110";
		Trees_din <= x"1a008d04";
		wait for Clk_period;
		Addr <=  "00001001001111";
		Trees_din <= x"001809e5";
		wait for Clk_period;
		Addr <=  "00001001010000";
		Trees_din <= x"ff6509e5";
		wait for Clk_period;
		Addr <=  "00001001010001";
		Trees_din <= x"02ff5708";
		wait for Clk_period;
		Addr <=  "00001001010010";
		Trees_din <= x"0b053004";
		wait for Clk_period;
		Addr <=  "00001001010011";
		Trees_din <= x"ff6c09e5";
		wait for Clk_period;
		Addr <=  "00001001010100";
		Trees_din <= x"ffef09e5";
		wait for Clk_period;
		Addr <=  "00001001010101";
		Trees_din <= x"1a00be08";
		wait for Clk_period;
		Addr <=  "00001001010110";
		Trees_din <= x"0efc2e04";
		wait for Clk_period;
		Addr <=  "00001001010111";
		Trees_din <= x"000e09e5";
		wait for Clk_period;
		Addr <=  "00001001011000";
		Trees_din <= x"ff7909e5";
		wait for Clk_period;
		Addr <=  "00001001011001";
		Trees_din <= x"1500a104";
		wait for Clk_period;
		Addr <=  "00001001011010";
		Trees_din <= x"009809e5";
		wait for Clk_period;
		Addr <=  "00001001011011";
		Trees_din <= x"ffb809e5";
		wait for Clk_period;
		Addr <=  "00001001011100";
		Trees_din <= x"040e6428";
		wait for Clk_period;
		Addr <=  "00001001011101";
		Trees_din <= x"03fb3a08";
		wait for Clk_period;
		Addr <=  "00001001011110";
		Trees_din <= x"01067004";
		wait for Clk_period;
		Addr <=  "00001001011111";
		Trees_din <= x"ffe309e5";
		wait for Clk_period;
		Addr <=  "00001001100000";
		Trees_din <= x"ff7709e5";
		wait for Clk_period;
		Addr <=  "00001001100001";
		Trees_din <= x"0d039d10";
		wait for Clk_period;
		Addr <=  "00001001100010";
		Trees_din <= x"10f75608";
		wait for Clk_period;
		Addr <=  "00001001100011";
		Trees_din <= x"0f002c04";
		wait for Clk_period;
		Addr <=  "00001001100100";
		Trees_din <= x"003009e5";
		wait for Clk_period;
		Addr <=  "00001001100101";
		Trees_din <= x"ff5c09e5";
		wait for Clk_period;
		Addr <=  "00001001100110";
		Trees_din <= x"18003c04";
		wait for Clk_period;
		Addr <=  "00001001100111";
		Trees_din <= x"005709e5";
		wait for Clk_period;
		Addr <=  "00001001101000";
		Trees_din <= x"000c09e5";
		wait for Clk_period;
		Addr <=  "00001001101001";
		Trees_din <= x"09005508";
		wait for Clk_period;
		Addr <=  "00001001101010";
		Trees_din <= x"13ffc104";
		wait for Clk_period;
		Addr <=  "00001001101011";
		Trees_din <= x"00d909e5";
		wait for Clk_period;
		Addr <=  "00001001101100";
		Trees_din <= x"000409e5";
		wait for Clk_period;
		Addr <=  "00001001101101";
		Trees_din <= x"1102c004";
		wait for Clk_period;
		Addr <=  "00001001101110";
		Trees_din <= x"ff7d09e5";
		wait for Clk_period;
		Addr <=  "00001001101111";
		Trees_din <= x"006c09e5";
		wait for Clk_period;
		Addr <=  "00001001110000";
		Trees_din <= x"030a7410";
		wait for Clk_period;
		Addr <=  "00001001110001";
		Trees_din <= x"16001e08";
		wait for Clk_period;
		Addr <=  "00001001110010";
		Trees_din <= x"0800ba04";
		wait for Clk_period;
		Addr <=  "00001001110011";
		Trees_din <= x"ffdd09e5";
		wait for Clk_period;
		Addr <=  "00001001110100";
		Trees_din <= x"006f09e5";
		wait for Clk_period;
		Addr <=  "00001001110101";
		Trees_din <= x"18003804";
		wait for Clk_period;
		Addr <=  "00001001110110";
		Trees_din <= x"000c09e5";
		wait for Clk_period;
		Addr <=  "00001001110111";
		Trees_din <= x"00bb09e5";
		wait for Clk_period;
		Addr <=  "00001001111000";
		Trees_din <= x"001209e5";
		wait for Clk_period;
		Addr <=  "00001001111001";
		Trees_din <= x"04041b34";
		wait for Clk_period;
		Addr <=  "00001001111010";
		Trees_din <= x"04fd5314";
		wait for Clk_period;
		Addr <=  "00001001111011";
		Trees_din <= x"0215a80c";
		wait for Clk_period;
		Addr <=  "00001001111100";
		Trees_din <= x"09003c08";
		wait for Clk_period;
		Addr <=  "00001001111101";
		Trees_din <= x"06f80d04";
		wait for Clk_period;
		Addr <=  "00001001111110";
		Trees_din <= x"ff9a0ad1";
		wait for Clk_period;
		Addr <=  "00001001111111";
		Trees_din <= x"00490ad1";
		wait for Clk_period;
		Addr <=  "00001010000000";
		Trees_din <= x"ff650ad1";
		wait for Clk_period;
		Addr <=  "00001010000001";
		Trees_din <= x"1a00bf04";
		wait for Clk_period;
		Addr <=  "00001010000010";
		Trees_din <= x"004a0ad1";
		wait for Clk_period;
		Addr <=  "00001010000011";
		Trees_din <= x"ffa70ad1";
		wait for Clk_period;
		Addr <=  "00001010000100";
		Trees_din <= x"06f5ff08";
		wait for Clk_period;
		Addr <=  "00001010000101";
		Trees_din <= x"1a008d04";
		wait for Clk_period;
		Addr <=  "00001010000110";
		Trees_din <= x"001a0ad1";
		wait for Clk_period;
		Addr <=  "00001010000111";
		Trees_din <= x"ff670ad1";
		wait for Clk_period;
		Addr <=  "00001010001000";
		Trees_din <= x"02ff5708";
		wait for Clk_period;
		Addr <=  "00001010001001";
		Trees_din <= x"04037804";
		wait for Clk_period;
		Addr <=  "00001010001010";
		Trees_din <= x"ff6f0ad1";
		wait for Clk_period;
		Addr <=  "00001010001011";
		Trees_din <= x"fff40ad1";
		wait for Clk_period;
		Addr <=  "00001010001100";
		Trees_din <= x"11013308";
		wait for Clk_period;
		Addr <=  "00001010001101";
		Trees_din <= x"02004a04";
		wait for Clk_period;
		Addr <=  "00001010001110";
		Trees_din <= x"003b0ad1";
		wait for Clk_period;
		Addr <=  "00001010001111";
		Trees_din <= x"ff780ad1";
		wait for Clk_period;
		Addr <=  "00001010010000";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00001010010001";
		Trees_din <= x"00750ad1";
		wait for Clk_period;
		Addr <=  "00001010010010";
		Trees_din <= x"ff860ad1";
		wait for Clk_period;
		Addr <=  "00001010010011";
		Trees_din <= x"040e6430";
		wait for Clk_period;
		Addr <=  "00001010010100";
		Trees_din <= x"07005a18";
		wait for Clk_period;
		Addr <=  "00001010010101";
		Trees_din <= x"0c03e210";
		wait for Clk_period;
		Addr <=  "00001010010110";
		Trees_din <= x"04065f08";
		wait for Clk_period;
		Addr <=  "00001010010111";
		Trees_din <= x"1701f304";
		wait for Clk_period;
		Addr <=  "00001010011000";
		Trees_din <= x"00180ad1";
		wait for Clk_period;
		Addr <=  "00001010011001";
		Trees_din <= x"ff650ad1";
		wait for Clk_period;
		Addr <=  "00001010011010";
		Trees_din <= x"0c03c404";
		wait for Clk_period;
		Addr <=  "00001010011011";
		Trees_din <= x"00390ad1";
		wait for Clk_period;
		Addr <=  "00001010011100";
		Trees_din <= x"ff560ad1";
		wait for Clk_period;
		Addr <=  "00001010011101";
		Trees_din <= x"1900a604";
		wait for Clk_period;
		Addr <=  "00001010011110";
		Trees_din <= x"00c70ad1";
		wait for Clk_period;
		Addr <=  "00001010011111";
		Trees_din <= x"001a0ad1";
		wait for Clk_period;
		Addr <=  "00001010100000";
		Trees_din <= x"0af7f108";
		wait for Clk_period;
		Addr <=  "00001010100001";
		Trees_din <= x"12009304";
		wait for Clk_period;
		Addr <=  "00001010100010";
		Trees_din <= x"ffe60ad1";
		wait for Clk_period;
		Addr <=  "00001010100011";
		Trees_din <= x"01000ad1";
		wait for Clk_period;
		Addr <=  "00001010100100";
		Trees_din <= x"17000208";
		wait for Clk_period;
		Addr <=  "00001010100101";
		Trees_din <= x"13f8ee04";
		wait for Clk_period;
		Addr <=  "00001010100110";
		Trees_din <= x"ff640ad1";
		wait for Clk_period;
		Addr <=  "00001010100111";
		Trees_din <= x"00230ad1";
		wait for Clk_period;
		Addr <=  "00001010101000";
		Trees_din <= x"19008204";
		wait for Clk_period;
		Addr <=  "00001010101001";
		Trees_din <= x"00110ad1";
		wait for Clk_period;
		Addr <=  "00001010101010";
		Trees_din <= x"ff560ad1";
		wait for Clk_period;
		Addr <=  "00001010101011";
		Trees_din <= x"030a7410";
		wait for Clk_period;
		Addr <=  "00001010101100";
		Trees_din <= x"16001e08";
		wait for Clk_period;
		Addr <=  "00001010101101";
		Trees_din <= x"00f9b904";
		wait for Clk_period;
		Addr <=  "00001010101110";
		Trees_din <= x"006a0ad1";
		wait for Clk_period;
		Addr <=  "00001010101111";
		Trees_din <= x"ffdb0ad1";
		wait for Clk_period;
		Addr <=  "00001010110000";
		Trees_din <= x"18003804";
		wait for Clk_period;
		Addr <=  "00001010110001";
		Trees_din <= x"00070ad1";
		wait for Clk_period;
		Addr <=  "00001010110010";
		Trees_din <= x"00b20ad1";
		wait for Clk_period;
		Addr <=  "00001010110011";
		Trees_din <= x"000f0ad1";
		wait for Clk_period;
		Addr <=  "00001010110100";
		Trees_din <= x"0401dd30";
		wait for Clk_period;
		Addr <=  "00001010110101";
		Trees_din <= x"03fbf60c";
		wait for Clk_period;
		Addr <=  "00001010110110";
		Trees_din <= x"0215a804";
		wait for Clk_period;
		Addr <=  "00001010110111";
		Trees_din <= x"ff660bbd";
		wait for Clk_period;
		Addr <=  "00001010111000";
		Trees_din <= x"0d01d904";
		wait for Clk_period;
		Addr <=  "00001010111001";
		Trees_din <= x"ffa90bbd";
		wait for Clk_period;
		Addr <=  "00001010111010";
		Trees_din <= x"00490bbd";
		wait for Clk_period;
		Addr <=  "00001010111011";
		Trees_din <= x"0c004308";
		wait for Clk_period;
		Addr <=  "00001010111100";
		Trees_din <= x"1b003604";
		wait for Clk_period;
		Addr <=  "00001010111101";
		Trees_din <= x"01020bbd";
		wait for Clk_period;
		Addr <=  "00001010111110";
		Trees_din <= x"ff970bbd";
		wait for Clk_period;
		Addr <=  "00001010111111";
		Trees_din <= x"0e045b10";
		wait for Clk_period;
		Addr <=  "00001011000000";
		Trees_din <= x"03fc2f08";
		wait for Clk_period;
		Addr <=  "00001011000001";
		Trees_din <= x"0d030704";
		wait for Clk_period;
		Addr <=  "00001011000010";
		Trees_din <= x"ffb00bbd";
		wait for Clk_period;
		Addr <=  "00001011000011";
		Trees_din <= x"00ce0bbd";
		wait for Clk_period;
		Addr <=  "00001011000100";
		Trees_din <= x"07004a04";
		wait for Clk_period;
		Addr <=  "00001011000101";
		Trees_din <= x"002e0bbd";
		wait for Clk_period;
		Addr <=  "00001011000110";
		Trees_din <= x"ff670bbd";
		wait for Clk_period;
		Addr <=  "00001011000111";
		Trees_din <= x"1a00e708";
		wait for Clk_period;
		Addr <=  "00001011001000";
		Trees_din <= x"00019004";
		wait for Clk_period;
		Addr <=  "00001011001001";
		Trees_din <= x"001d0bbd";
		wait for Clk_period;
		Addr <=  "00001011001010";
		Trees_din <= x"ff9e0bbd";
		wait for Clk_period;
		Addr <=  "00001011001011";
		Trees_din <= x"00d30bbd";
		wait for Clk_period;
		Addr <=  "00001011001100";
		Trees_din <= x"04065f1c";
		wait for Clk_period;
		Addr <=  "00001011001101";
		Trees_din <= x"06f4ea08";
		wait for Clk_period;
		Addr <=  "00001011001110";
		Trees_din <= x"0e040704";
		wait for Clk_period;
		Addr <=  "00001011001111";
		Trees_din <= x"ff670bbd";
		wait for Clk_period;
		Addr <=  "00001011010000";
		Trees_din <= x"007c0bbd";
		wait for Clk_period;
		Addr <=  "00001011010001";
		Trees_din <= x"1702c810";
		wait for Clk_period;
		Addr <=  "00001011010010";
		Trees_din <= x"1601bb08";
		wait for Clk_period;
		Addr <=  "00001011010011";
		Trees_din <= x"02007704";
		wait for Clk_period;
		Addr <=  "00001011010100";
		Trees_din <= x"ff960bbd";
		wait for Clk_period;
		Addr <=  "00001011010101";
		Trees_din <= x"002e0bbd";
		wait for Clk_period;
		Addr <=  "00001011010110";
		Trees_din <= x"07005104";
		wait for Clk_period;
		Addr <=  "00001011010111";
		Trees_din <= x"ffa70bbd";
		wait for Clk_period;
		Addr <=  "00001011011000";
		Trees_din <= x"007e0bbd";
		wait for Clk_period;
		Addr <=  "00001011011001";
		Trees_din <= x"ff700bbd";
		wait for Clk_period;
		Addr <=  "00001011011010";
		Trees_din <= x"040e641c";
		wait for Clk_period;
		Addr <=  "00001011011011";
		Trees_din <= x"1600010c";
		wait for Clk_period;
		Addr <=  "00001011011100";
		Trees_din <= x"0d005808";
		wait for Clk_period;
		Addr <=  "00001011011101";
		Trees_din <= x"16000004";
		wait for Clk_period;
		Addr <=  "00001011011110";
		Trees_din <= x"003b0bbd";
		wait for Clk_period;
		Addr <=  "00001011011111";
		Trees_din <= x"00ed0bbd";
		wait for Clk_period;
		Addr <=  "00001011100000";
		Trees_din <= x"ffe60bbd";
		wait for Clk_period;
		Addr <=  "00001011100001";
		Trees_din <= x"07005a08";
		wait for Clk_period;
		Addr <=  "00001011100010";
		Trees_din <= x"01036504";
		wait for Clk_period;
		Addr <=  "00001011100011";
		Trees_din <= x"004a0bbd";
		wait for Clk_period;
		Addr <=  "00001011100100";
		Trees_din <= x"fffe0bbd";
		wait for Clk_period;
		Addr <=  "00001011100101";
		Trees_din <= x"18004a04";
		wait for Clk_period;
		Addr <=  "00001011100110";
		Trees_din <= x"ff940bbd";
		wait for Clk_period;
		Addr <=  "00001011100111";
		Trees_din <= x"00650bbd";
		wait for Clk_period;
		Addr <=  "00001011101000";
		Trees_din <= x"030a740c";
		wait for Clk_period;
		Addr <=  "00001011101001";
		Trees_din <= x"08000904";
		wait for Clk_period;
		Addr <=  "00001011101010";
		Trees_din <= x"000f0bbd";
		wait for Clk_period;
		Addr <=  "00001011101011";
		Trees_din <= x"16001e04";
		wait for Clk_period;
		Addr <=  "00001011101100";
		Trees_din <= x"00290bbd";
		wait for Clk_period;
		Addr <=  "00001011101101";
		Trees_din <= x"00a90bbd";
		wait for Clk_period;
		Addr <=  "00001011101110";
		Trees_din <= x"000b0bbd";
		wait for Clk_period;
		Addr <=  "00001011101111";
		Trees_din <= x"0401dd2c";
		wait for Clk_period;
		Addr <=  "00001011110000";
		Trees_din <= x"03fbf608";
		wait for Clk_period;
		Addr <=  "00001011110001";
		Trees_din <= x"0215a804";
		wait for Clk_period;
		Addr <=  "00001011110010";
		Trees_din <= x"ff660ca1";
		wait for Clk_period;
		Addr <=  "00001011110011";
		Trees_din <= x"ffff0ca1";
		wait for Clk_period;
		Addr <=  "00001011110100";
		Trees_din <= x"0c004308";
		wait for Clk_period;
		Addr <=  "00001011110101";
		Trees_din <= x"1b003604";
		wait for Clk_period;
		Addr <=  "00001011110110";
		Trees_din <= x"00d20ca1";
		wait for Clk_period;
		Addr <=  "00001011110111";
		Trees_din <= x"ff9c0ca1";
		wait for Clk_period;
		Addr <=  "00001011111000";
		Trees_din <= x"0e045b10";
		wait for Clk_period;
		Addr <=  "00001011111001";
		Trees_din <= x"03fc2f08";
		wait for Clk_period;
		Addr <=  "00001011111010";
		Trees_din <= x"10046604";
		wait for Clk_period;
		Addr <=  "00001011111011";
		Trees_din <= x"ffad0ca1";
		wait for Clk_period;
		Addr <=  "00001011111100";
		Trees_din <= x"00ce0ca1";
		wait for Clk_period;
		Addr <=  "00001011111101";
		Trees_din <= x"07004a04";
		wait for Clk_period;
		Addr <=  "00001011111110";
		Trees_din <= x"002c0ca1";
		wait for Clk_period;
		Addr <=  "00001011111111";
		Trees_din <= x"ff680ca1";
		wait for Clk_period;
		Addr <=  "00001100000000";
		Trees_din <= x"0bfb0108";
		wait for Clk_period;
		Addr <=  "00001100000001";
		Trees_din <= x"1601ee04";
		wait for Clk_period;
		Addr <=  "00001100000010";
		Trees_din <= x"00140ca1";
		wait for Clk_period;
		Addr <=  "00001100000011";
		Trees_din <= x"00cc0ca1";
		wait for Clk_period;
		Addr <=  "00001100000100";
		Trees_din <= x"ffa30ca1";
		wait for Clk_period;
		Addr <=  "00001100000101";
		Trees_din <= x"04065f18";
		wait for Clk_period;
		Addr <=  "00001100000110";
		Trees_din <= x"06f4ea08";
		wait for Clk_period;
		Addr <=  "00001100000111";
		Trees_din <= x"0e040704";
		wait for Clk_period;
		Addr <=  "00001100001000";
		Trees_din <= x"ff6a0ca1";
		wait for Clk_period;
		Addr <=  "00001100001001";
		Trees_din <= x"00690ca1";
		wait for Clk_period;
		Addr <=  "00001100001010";
		Trees_din <= x"1702c80c";
		wait for Clk_period;
		Addr <=  "00001100001011";
		Trees_din <= x"12fed404";
		wait for Clk_period;
		Addr <=  "00001100001100";
		Trees_din <= x"ff7a0ca1";
		wait for Clk_period;
		Addr <=  "00001100001101";
		Trees_din <= x"1b002c04";
		wait for Clk_period;
		Addr <=  "00001100001110";
		Trees_din <= x"ff910ca1";
		wait for Clk_period;
		Addr <=  "00001100001111";
		Trees_din <= x"00420ca1";
		wait for Clk_period;
		Addr <=  "00001100010000";
		Trees_din <= x"ff740ca1";
		wait for Clk_period;
		Addr <=  "00001100010001";
		Trees_din <= x"040e6420";
		wait for Clk_period;
		Addr <=  "00001100010010";
		Trees_din <= x"15009f10";
		wait for Clk_period;
		Addr <=  "00001100010011";
		Trees_din <= x"0d033b08";
		wait for Clk_period;
		Addr <=  "00001100010100";
		Trees_din <= x"16011904";
		wait for Clk_period;
		Addr <=  "00001100010101";
		Trees_din <= x"002e0ca1";
		wait for Clk_period;
		Addr <=  "00001100010110";
		Trees_din <= x"ffc20ca1";
		wait for Clk_period;
		Addr <=  "00001100010111";
		Trees_din <= x"0c024504";
		wait for Clk_period;
		Addr <=  "00001100011000";
		Trees_din <= x"00990ca1";
		wait for Clk_period;
		Addr <=  "00001100011001";
		Trees_din <= x"000a0ca1";
		wait for Clk_period;
		Addr <=  "00001100011010";
		Trees_din <= x"1c002508";
		wait for Clk_period;
		Addr <=  "00001100011011";
		Trees_din <= x"0b046404";
		wait for Clk_period;
		Addr <=  "00001100011100";
		Trees_din <= x"ff700ca1";
		wait for Clk_period;
		Addr <=  "00001100011101";
		Trees_din <= x"00620ca1";
		wait for Clk_period;
		Addr <=  "00001100011110";
		Trees_din <= x"05f8b404";
		wait for Clk_period;
		Addr <=  "00001100011111";
		Trees_din <= x"ff880ca1";
		wait for Clk_period;
		Addr <=  "00001100100000";
		Trees_din <= x"007d0ca1";
		wait for Clk_period;
		Addr <=  "00001100100001";
		Trees_din <= x"12fbf704";
		wait for Clk_period;
		Addr <=  "00001100100010";
		Trees_din <= x"fff60ca1";
		wait for Clk_period;
		Addr <=  "00001100100011";
		Trees_din <= x"05f8f708";
		wait for Clk_period;
		Addr <=  "00001100100100";
		Trees_din <= x"0bf96504";
		wait for Clk_period;
		Addr <=  "00001100100101";
		Trees_din <= x"ffbe0ca1";
		wait for Clk_period;
		Addr <=  "00001100100110";
		Trees_din <= x"00680ca1";
		wait for Clk_period;
		Addr <=  "00001100100111";
		Trees_din <= x"00a20ca1";
		wait for Clk_period;
		Addr <=  "00001100101000";
		Trees_din <= x"0401dd24";
		wait for Clk_period;
		Addr <=  "00001100101001";
		Trees_din <= x"03fbf608";
		wait for Clk_period;
		Addr <=  "00001100101010";
		Trees_din <= x"0215a804";
		wait for Clk_period;
		Addr <=  "00001100101011";
		Trees_din <= x"ff670d85";
		wait for Clk_period;
		Addr <=  "00001100101100";
		Trees_din <= x"00050d85";
		wait for Clk_period;
		Addr <=  "00001100101101";
		Trees_din <= x"0c004308";
		wait for Clk_period;
		Addr <=  "00001100101110";
		Trees_din <= x"1b003604";
		wait for Clk_period;
		Addr <=  "00001100101111";
		Trees_din <= x"00b70d85";
		wait for Clk_period;
		Addr <=  "00001100110000";
		Trees_din <= x"ffa10d85";
		wait for Clk_period;
		Addr <=  "00001100110001";
		Trees_din <= x"1103a608";
		wait for Clk_period;
		Addr <=  "00001100110010";
		Trees_din <= x"03fc2f04";
		wait for Clk_period;
		Addr <=  "00001100110011";
		Trees_din <= x"00530d85";
		wait for Clk_period;
		Addr <=  "00001100110100";
		Trees_din <= x"ff6a0d85";
		wait for Clk_period;
		Addr <=  "00001100110101";
		Trees_din <= x"12034508";
		wait for Clk_period;
		Addr <=  "00001100110110";
		Trees_din <= x"1a00d904";
		wait for Clk_period;
		Addr <=  "00001100110111";
		Trees_din <= x"ffff0d85";
		wait for Clk_period;
		Addr <=  "00001100111000";
		Trees_din <= x"01300d85";
		wait for Clk_period;
		Addr <=  "00001100111001";
		Trees_din <= x"ff860d85";
		wait for Clk_period;
		Addr <=  "00001100111010";
		Trees_din <= x"040a4a28";
		wait for Clk_period;
		Addr <=  "00001100111011";
		Trees_din <= x"1d003608";
		wait for Clk_period;
		Addr <=  "00001100111100";
		Trees_din <= x"11006c04";
		wait for Clk_period;
		Addr <=  "00001100111101";
		Trees_din <= x"002d0d85";
		wait for Clk_period;
		Addr <=  "00001100111110";
		Trees_din <= x"ff5f0d85";
		wait for Clk_period;
		Addr <=  "00001100111111";
		Trees_din <= x"1c002c10";
		wait for Clk_period;
		Addr <=  "00001101000000";
		Trees_din <= x"0801fa08";
		wait for Clk_period;
		Addr <=  "00001101000001";
		Trees_din <= x"00fd6404";
		wait for Clk_period;
		Addr <=  "00001101000010";
		Trees_din <= x"00010d85";
		wait for Clk_period;
		Addr <=  "00001101000011";
		Trees_din <= x"00a10d85";
		wait for Clk_period;
		Addr <=  "00001101000100";
		Trees_din <= x"1400f204";
		wait for Clk_period;
		Addr <=  "00001101000101";
		Trees_din <= x"00660d85";
		wait for Clk_period;
		Addr <=  "00001101000110";
		Trees_din <= x"ff950d85";
		wait for Clk_period;
		Addr <=  "00001101000111";
		Trees_din <= x"16000508";
		wait for Clk_period;
		Addr <=  "00001101001000";
		Trees_din <= x"0e020804";
		wait for Clk_period;
		Addr <=  "00001101001001";
		Trees_din <= x"00910d85";
		wait for Clk_period;
		Addr <=  "00001101001010";
		Trees_din <= x"ff7f0d85";
		wait for Clk_period;
		Addr <=  "00001101001011";
		Trees_din <= x"00fce804";
		wait for Clk_period;
		Addr <=  "00001101001100";
		Trees_din <= x"002d0d85";
		wait for Clk_period;
		Addr <=  "00001101001101";
		Trees_din <= x"ffd30d85";
		wait for Clk_period;
		Addr <=  "00001101001110";
		Trees_din <= x"07005510";
		wait for Clk_period;
		Addr <=  "00001101001111";
		Trees_din <= x"0bf98b04";
		wait for Clk_period;
		Addr <=  "00001101010000";
		Trees_din <= x"ffb30d85";
		wait for Clk_period;
		Addr <=  "00001101010001";
		Trees_din <= x"030a7408";
		wait for Clk_period;
		Addr <=  "00001101010010";
		Trees_din <= x"08035604";
		wait for Clk_period;
		Addr <=  "00001101010011";
		Trees_din <= x"00b60d85";
		wait for Clk_period;
		Addr <=  "00001101010100";
		Trees_din <= x"00300d85";
		wait for Clk_period;
		Addr <=  "00001101010101";
		Trees_din <= x"fffc0d85";
		wait for Clk_period;
		Addr <=  "00001101010110";
		Trees_din <= x"13f88908";
		wait for Clk_period;
		Addr <=  "00001101010111";
		Trees_din <= x"13f83104";
		wait for Clk_period;
		Addr <=  "00001101011000";
		Trees_din <= x"002e0d85";
		wait for Clk_period;
		Addr <=  "00001101011001";
		Trees_din <= x"ff560d85";
		wait for Clk_period;
		Addr <=  "00001101011010";
		Trees_din <= x"1e007008";
		wait for Clk_period;
		Addr <=  "00001101011011";
		Trees_din <= x"18004204";
		wait for Clk_period;
		Addr <=  "00001101011100";
		Trees_din <= x"002e0d85";
		wait for Clk_period;
		Addr <=  "00001101011101";
		Trees_din <= x"ff510d85";
		wait for Clk_period;
		Addr <=  "00001101011110";
		Trees_din <= x"02fba504";
		wait for Clk_period;
		Addr <=  "00001101011111";
		Trees_din <= x"ffb70d85";
		wait for Clk_period;
		Addr <=  "00001101100000";
		Trees_din <= x"007f0d85";
		wait for Clk_period;
		Addr <=  "00001101100001";
		Trees_din <= x"0401dd24";
		wait for Clk_period;
		Addr <=  "00001101100010";
		Trees_din <= x"03fbf608";
		wait for Clk_period;
		Addr <=  "00001101100011";
		Trees_din <= x"0215a804";
		wait for Clk_period;
		Addr <=  "00001101100100";
		Trees_din <= x"ff680e39";
		wait for Clk_period;
		Addr <=  "00001101100101";
		Trees_din <= x"00100e39";
		wait for Clk_period;
		Addr <=  "00001101100110";
		Trees_din <= x"0c004308";
		wait for Clk_period;
		Addr <=  "00001101100111";
		Trees_din <= x"1b003604";
		wait for Clk_period;
		Addr <=  "00001101101000";
		Trees_din <= x"00a40e39";
		wait for Clk_period;
		Addr <=  "00001101101001";
		Trees_din <= x"ffa60e39";
		wait for Clk_period;
		Addr <=  "00001101101010";
		Trees_din <= x"1103a608";
		wait for Clk_period;
		Addr <=  "00001101101011";
		Trees_din <= x"03fc2f04";
		wait for Clk_period;
		Addr <=  "00001101101100";
		Trees_din <= x"004c0e39";
		wait for Clk_period;
		Addr <=  "00001101101101";
		Trees_din <= x"ff6c0e39";
		wait for Clk_period;
		Addr <=  "00001101101110";
		Trees_din <= x"12034508";
		wait for Clk_period;
		Addr <=  "00001101101111";
		Trees_din <= x"1a00d904";
		wait for Clk_period;
		Addr <=  "00001101110000";
		Trees_din <= x"fffd0e39";
		wait for Clk_period;
		Addr <=  "00001101110001";
		Trees_din <= x"00fe0e39";
		wait for Clk_period;
		Addr <=  "00001101110010";
		Trees_din <= x"ff8b0e39";
		wait for Clk_period;
		Addr <=  "00001101110011";
		Trees_din <= x"040e6424";
		wait for Clk_period;
		Addr <=  "00001101110100";
		Trees_din <= x"03fb1e04";
		wait for Clk_period;
		Addr <=  "00001101110101";
		Trees_din <= x"ff860e39";
		wait for Clk_period;
		Addr <=  "00001101110110";
		Trees_din <= x"07005a10";
		wait for Clk_period;
		Addr <=  "00001101110111";
		Trees_din <= x"07005008";
		wait for Clk_period;
		Addr <=  "00001101111000";
		Trees_din <= x"040c1204";
		wait for Clk_period;
		Addr <=  "00001101111001";
		Trees_din <= x"ffb40e39";
		wait for Clk_period;
		Addr <=  "00001101111010";
		Trees_din <= x"007a0e39";
		wait for Clk_period;
		Addr <=  "00001101111011";
		Trees_din <= x"06f4a504";
		wait for Clk_period;
		Addr <=  "00001101111100";
		Trees_din <= x"fff60e39";
		wait for Clk_period;
		Addr <=  "00001101111101";
		Trees_din <= x"00340e39";
		wait for Clk_period;
		Addr <=  "00001101111110";
		Trees_din <= x"0af7f108";
		wait for Clk_period;
		Addr <=  "00001101111111";
		Trees_din <= x"1a00b104";
		wait for Clk_period;
		Addr <=  "00001110000000";
		Trees_din <= x"00c10e39";
		wait for Clk_period;
		Addr <=  "00001110000001";
		Trees_din <= x"ffe50e39";
		wait for Clk_period;
		Addr <=  "00001110000010";
		Trees_din <= x"17000204";
		wait for Clk_period;
		Addr <=  "00001110000011";
		Trees_din <= x"fff20e39";
		wait for Clk_period;
		Addr <=  "00001110000100";
		Trees_din <= x"ff720e39";
		wait for Clk_period;
		Addr <=  "00001110000101";
		Trees_din <= x"05f95310";
		wait for Clk_period;
		Addr <=  "00001110000110";
		Trees_din <= x"0f00b308";
		wait for Clk_period;
		Addr <=  "00001110000111";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00001110001000";
		Trees_din <= x"00850e39";
		wait for Clk_period;
		Addr <=  "00001110001001";
		Trees_din <= x"00230e39";
		wait for Clk_period;
		Addr <=  "00001110001010";
		Trees_din <= x"0e01ff04";
		wait for Clk_period;
		Addr <=  "00001110001011";
		Trees_din <= x"00130e39";
		wait for Clk_period;
		Addr <=  "00001110001100";
		Trees_din <= x"ff8d0e39";
		wait for Clk_period;
		Addr <=  "00001110001101";
		Trees_din <= x"00940e39";
		wait for Clk_period;
		Addr <=  "00001110001110";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00001110001111";
		Trees_din <= x"0401dd2c";
		wait for Clk_period;
		Addr <=  "00001110010000";
		Trees_din <= x"03fbf608";
		wait for Clk_period;
		Addr <=  "00001110010001";
		Trees_din <= x"0215a804";
		wait for Clk_period;
		Addr <=  "00001110010010";
		Trees_din <= x"ff680f29";
		wait for Clk_period;
		Addr <=  "00001110010011";
		Trees_din <= x"00160f29";
		wait for Clk_period;
		Addr <=  "00001110010100";
		Trees_din <= x"05fe7018";
		wait for Clk_period;
		Addr <=  "00001110010101";
		Trees_din <= x"0e045b0c";
		wait for Clk_period;
		Addr <=  "00001110010110";
		Trees_din <= x"1c002304";
		wait for Clk_period;
		Addr <=  "00001110010111";
		Trees_din <= x"002a0f29";
		wait for Clk_period;
		Addr <=  "00001110011000";
		Trees_din <= x"0f03fb04";
		wait for Clk_period;
		Addr <=  "00001110011001";
		Trees_din <= x"ff6e0f29";
		wait for Clk_period;
		Addr <=  "00001110011010";
		Trees_din <= x"000e0f29";
		wait for Clk_period;
		Addr <=  "00001110011011";
		Trees_din <= x"20040008";
		wait for Clk_period;
		Addr <=  "00001110011100";
		Trees_din <= x"1a00e504";
		wait for Clk_period;
		Addr <=  "00001110011101";
		Trees_din <= x"000d0f29";
		wait for Clk_period;
		Addr <=  "00001110011110";
		Trees_din <= x"008f0f29";
		wait for Clk_period;
		Addr <=  "00001110011111";
		Trees_din <= x"ffac0f29";
		wait for Clk_period;
		Addr <=  "00001110100000";
		Trees_din <= x"05fefa04";
		wait for Clk_period;
		Addr <=  "00001110100001";
		Trees_din <= x"00fa0f29";
		wait for Clk_period;
		Addr <=  "00001110100010";
		Trees_din <= x"1402e804";
		wait for Clk_period;
		Addr <=  "00001110100011";
		Trees_din <= x"ff8c0f29";
		wait for Clk_period;
		Addr <=  "00001110100100";
		Trees_din <= x"00130f29";
		wait for Clk_period;
		Addr <=  "00001110100101";
		Trees_din <= x"04065f20";
		wait for Clk_period;
		Addr <=  "00001110100110";
		Trees_din <= x"1701f318";
		wait for Clk_period;
		Addr <=  "00001110100111";
		Trees_din <= x"0e01ba0c";
		wait for Clk_period;
		Addr <=  "00001110101000";
		Trees_din <= x"1a008d04";
		wait for Clk_period;
		Addr <=  "00001110101001";
		Trees_din <= x"008b0f29";
		wait for Clk_period;
		Addr <=  "00001110101010";
		Trees_din <= x"17003704";
		wait for Clk_period;
		Addr <=  "00001110101011";
		Trees_din <= x"ff8f0f29";
		wait for Clk_period;
		Addr <=  "00001110101100";
		Trees_din <= x"00170f29";
		wait for Clk_period;
		Addr <=  "00001110101101";
		Trees_din <= x"1900a908";
		wait for Clk_period;
		Addr <=  "00001110101110";
		Trees_din <= x"07005604";
		wait for Clk_period;
		Addr <=  "00001110101111";
		Trees_din <= x"00d30f29";
		wait for Clk_period;
		Addr <=  "00001110110000";
		Trees_din <= x"000e0f29";
		wait for Clk_period;
		Addr <=  "00001110110001";
		Trees_din <= x"ff850f29";
		wait for Clk_period;
		Addr <=  "00001110110010";
		Trees_din <= x"0c018c04";
		wait for Clk_period;
		Addr <=  "00001110110011";
		Trees_din <= x"ff6b0f29";
		wait for Clk_period;
		Addr <=  "00001110110100";
		Trees_din <= x"00120f29";
		wait for Clk_period;
		Addr <=  "00001110110101";
		Trees_din <= x"10028414";
		wait for Clk_period;
		Addr <=  "00001110110110";
		Trees_din <= x"1a008b04";
		wait for Clk_period;
		Addr <=  "00001110110111";
		Trees_din <= x"00b40f29";
		wait for Clk_period;
		Addr <=  "00001110111000";
		Trees_din <= x"1500a008";
		wait for Clk_period;
		Addr <=  "00001110111001";
		Trees_din <= x"1e006304";
		wait for Clk_period;
		Addr <=  "00001110111010";
		Trees_din <= x"ff5b0f29";
		wait for Clk_period;
		Addr <=  "00001110111011";
		Trees_din <= x"fff20f29";
		wait for Clk_period;
		Addr <=  "00001110111100";
		Trees_din <= x"0202d904";
		wait for Clk_period;
		Addr <=  "00001110111101";
		Trees_din <= x"00560f29";
		wait for Clk_period;
		Addr <=  "00001110111110";
		Trees_din <= x"ff7f0f29";
		wait for Clk_period;
		Addr <=  "00001110111111";
		Trees_din <= x"18005210";
		wait for Clk_period;
		Addr <=  "00001111000000";
		Trees_din <= x"1f000008";
		wait for Clk_period;
		Addr <=  "00001111000001";
		Trees_din <= x"0e024b04";
		wait for Clk_period;
		Addr <=  "00001111000010";
		Trees_din <= x"005b0f29";
		wait for Clk_period;
		Addr <=  "00001111000011";
		Trees_din <= x"ffc80f29";
		wait for Clk_period;
		Addr <=  "00001111000100";
		Trees_din <= x"12fe8304";
		wait for Clk_period;
		Addr <=  "00001111000101";
		Trees_din <= x"00410f29";
		wait for Clk_period;
		Addr <=  "00001111000110";
		Trees_din <= x"ff590f29";
		wait for Clk_period;
		Addr <=  "00001111000111";
		Trees_din <= x"14007804";
		wait for Clk_period;
		Addr <=  "00001111001000";
		Trees_din <= x"ffe60f29";
		wait for Clk_period;
		Addr <=  "00001111001001";
		Trees_din <= x"ff810f29";
		wait for Clk_period;
		Addr <=  "00001111001010";
		Trees_din <= x"04007b1c";
		wait for Clk_period;
		Addr <=  "00001111001011";
		Trees_din <= x"03fc1508";
		wait for Clk_period;
		Addr <=  "00001111001100";
		Trees_din <= x"1c005004";
		wait for Clk_period;
		Addr <=  "00001111001101";
		Trees_din <= x"ff690fed";
		wait for Clk_period;
		Addr <=  "00001111001110";
		Trees_din <= x"002c0fed";
		wait for Clk_period;
		Addr <=  "00001111001111";
		Trees_din <= x"0afce410";
		wait for Clk_period;
		Addr <=  "00001111010000";
		Trees_din <= x"12011308";
		wait for Clk_period;
		Addr <=  "00001111010001";
		Trees_din <= x"1a00d104";
		wait for Clk_period;
		Addr <=  "00001111010010";
		Trees_din <= x"ffac0fed";
		wait for Clk_period;
		Addr <=  "00001111010011";
		Trees_din <= x"01090fed";
		wait for Clk_period;
		Addr <=  "00001111010100";
		Trees_din <= x"0f02c604";
		wait for Clk_period;
		Addr <=  "00001111010101";
		Trees_din <= x"ff7e0fed";
		wait for Clk_period;
		Addr <=  "00001111010110";
		Trees_din <= x"00360fed";
		wait for Clk_period;
		Addr <=  "00001111010111";
		Trees_din <= x"ff760fed";
		wait for Clk_period;
		Addr <=  "00001111011000";
		Trees_din <= x"0404aa18";
		wait for Clk_period;
		Addr <=  "00001111011001";
		Trees_din <= x"02ff8608";
		wait for Clk_period;
		Addr <=  "00001111011010";
		Trees_din <= x"0b053004";
		wait for Clk_period;
		Addr <=  "00001111011011";
		Trees_din <= x"ff6f0fed";
		wait for Clk_period;
		Addr <=  "00001111011100";
		Trees_din <= x"00030fed";
		wait for Clk_period;
		Addr <=  "00001111011101";
		Trees_din <= x"06f4ea04";
		wait for Clk_period;
		Addr <=  "00001111011110";
		Trees_din <= x"ff7b0fed";
		wait for Clk_period;
		Addr <=  "00001111011111";
		Trees_din <= x"07005204";
		wait for Clk_period;
		Addr <=  "00001111100000";
		Trees_din <= x"ff960fed";
		wait for Clk_period;
		Addr <=  "00001111100001";
		Trees_din <= x"0b04c104";
		wait for Clk_period;
		Addr <=  "00001111100010";
		Trees_din <= x"00580fed";
		wait for Clk_period;
		Addr <=  "00001111100011";
		Trees_din <= x"ff990fed";
		wait for Clk_period;
		Addr <=  "00001111100100";
		Trees_din <= x"0d03ab1c";
		wait for Clk_period;
		Addr <=  "00001111100101";
		Trees_din <= x"1600010c";
		wait for Clk_period;
		Addr <=  "00001111100110";
		Trees_din <= x"00fba504";
		wait for Clk_period;
		Addr <=  "00001111100111";
		Trees_din <= x"ffec0fed";
		wait for Clk_period;
		Addr <=  "00001111101000";
		Trees_din <= x"1003b904";
		wait for Clk_period;
		Addr <=  "00001111101001";
		Trees_din <= x"00b70fed";
		wait for Clk_period;
		Addr <=  "00001111101010";
		Trees_din <= x"001f0fed";
		wait for Clk_period;
		Addr <=  "00001111101011";
		Trees_din <= x"07005808";
		wait for Clk_period;
		Addr <=  "00001111101100";
		Trees_din <= x"1900a804";
		wait for Clk_period;
		Addr <=  "00001111101101";
		Trees_din <= x"002b0fed";
		wait for Clk_period;
		Addr <=  "00001111101110";
		Trees_din <= x"ffde0fed";
		wait for Clk_period;
		Addr <=  "00001111101111";
		Trees_din <= x"1104d504";
		wait for Clk_period;
		Addr <=  "00001111110000";
		Trees_din <= x"ffd40fed";
		wait for Clk_period;
		Addr <=  "00001111110001";
		Trees_din <= x"00bd0fed";
		wait for Clk_period;
		Addr <=  "00001111110010";
		Trees_din <= x"0900550c";
		wait for Clk_period;
		Addr <=  "00001111110011";
		Trees_din <= x"01fbcc04";
		wait for Clk_period;
		Addr <=  "00001111110100";
		Trees_din <= x"00020fed";
		wait for Clk_period;
		Addr <=  "00001111110101";
		Trees_din <= x"06f37104";
		wait for Clk_period;
		Addr <=  "00001111110110";
		Trees_din <= x"003c0fed";
		wait for Clk_period;
		Addr <=  "00001111110111";
		Trees_din <= x"00c60fed";
		wait for Clk_period;
		Addr <=  "00001111111000";
		Trees_din <= x"17002c04";
		wait for Clk_period;
		Addr <=  "00001111111001";
		Trees_din <= x"00080fed";
		wait for Clk_period;
		Addr <=  "00001111111010";
		Trees_din <= x"ffaa0fed";
		wait for Clk_period;
		Addr <=  "00001111111011";
		Trees_din <= x"03fb1e0c";
		wait for Clk_period;
		Addr <=  "00001111111100";
		Trees_din <= x"0215a808";
		wait for Clk_period;
		Addr <=  "00001111111101";
		Trees_din <= x"00ff7304";
		wait for Clk_period;
		Addr <=  "00001111111110";
		Trees_din <= x"fff510b1";
		wait for Clk_period;
		Addr <=  "00001111111111";
		Trees_din <= x"ff6910b1";
		wait for Clk_period;
		Addr <=  "00010000000000";
		Trees_din <= x"003710b1";
		wait for Clk_period;
		Addr <=  "00010000000001";
		Trees_din <= x"0404aa28";
		wait for Clk_period;
		Addr <=  "00010000000010";
		Trees_din <= x"01fdac10";
		wait for Clk_period;
		Addr <=  "00010000000011";
		Trees_din <= x"0307f50c";
		wait for Clk_period;
		Addr <=  "00010000000100";
		Trees_din <= x"0d02e908";
		wait for Clk_period;
		Addr <=  "00010000000101";
		Trees_din <= x"0afb0304";
		wait for Clk_period;
		Addr <=  "00010000000110";
		Trees_din <= x"00f810b1";
		wait for Clk_period;
		Addr <=  "00010000000111";
		Trees_din <= x"001510b1";
		wait for Clk_period;
		Addr <=  "00010000001000";
		Trees_din <= x"ff9e10b1";
		wait for Clk_period;
		Addr <=  "00010000001001";
		Trees_din <= x"ff8c10b1";
		wait for Clk_period;
		Addr <=  "00010000001010";
		Trees_din <= x"1602f310";
		wait for Clk_period;
		Addr <=  "00010000001011";
		Trees_din <= x"01056508";
		wait for Clk_period;
		Addr <=  "00010000001100";
		Trees_din <= x"17009e04";
		wait for Clk_period;
		Addr <=  "00010000001101";
		Trees_din <= x"ff7d10b1";
		wait for Clk_period;
		Addr <=  "00010000001110";
		Trees_din <= x"001910b1";
		wait for Clk_period;
		Addr <=  "00010000001111";
		Trees_din <= x"06f51304";
		wait for Clk_period;
		Addr <=  "00010000010000";
		Trees_din <= x"ff8f10b1";
		wait for Clk_period;
		Addr <=  "00010000010001";
		Trees_din <= x"005810b1";
		wait for Clk_period;
		Addr <=  "00010000010010";
		Trees_din <= x"0308a904";
		wait for Clk_period;
		Addr <=  "00010000010011";
		Trees_din <= x"ff6b10b1";
		wait for Clk_period;
		Addr <=  "00010000010100";
		Trees_din <= x"001e10b1";
		wait for Clk_period;
		Addr <=  "00010000010101";
		Trees_din <= x"0d039d18";
		wait for Clk_period;
		Addr <=  "00010000010110";
		Trees_din <= x"02091310";
		wait for Clk_period;
		Addr <=  "00010000010111";
		Trees_din <= x"0b04f208";
		wait for Clk_period;
		Addr <=  "00010000011000";
		Trees_din <= x"05fcbb04";
		wait for Clk_period;
		Addr <=  "00010000011001";
		Trees_din <= x"ffe210b1";
		wait for Clk_period;
		Addr <=  "00010000011010";
		Trees_din <= x"001d10b1";
		wait for Clk_period;
		Addr <=  "00010000011011";
		Trees_din <= x"19009e04";
		wait for Clk_period;
		Addr <=  "00010000011100";
		Trees_din <= x"fff810b1";
		wait for Clk_period;
		Addr <=  "00010000011101";
		Trees_din <= x"00b110b1";
		wait for Clk_period;
		Addr <=  "00010000011110";
		Trees_din <= x"0afccf04";
		wait for Clk_period;
		Addr <=  "00010000011111";
		Trees_din <= x"00f010b1";
		wait for Clk_period;
		Addr <=  "00010000100000";
		Trees_din <= x"fff910b1";
		wait for Clk_period;
		Addr <=  "00010000100001";
		Trees_din <= x"0900560c";
		wait for Clk_period;
		Addr <=  "00010000100010";
		Trees_din <= x"04094204";
		wait for Clk_period;
		Addr <=  "00010000100011";
		Trees_din <= x"00ab10b1";
		wait for Clk_period;
		Addr <=  "00010000100100";
		Trees_din <= x"05fb8404";
		wait for Clk_period;
		Addr <=  "00010000100101";
		Trees_din <= x"005f10b1";
		wait for Clk_period;
		Addr <=  "00010000100110";
		Trees_din <= x"ffb110b1";
		wait for Clk_period;
		Addr <=  "00010000100111";
		Trees_din <= x"06f57808";
		wait for Clk_period;
		Addr <=  "00010000101000";
		Trees_din <= x"12021e04";
		wait for Clk_period;
		Addr <=  "00010000101001";
		Trees_din <= x"fffc10b1";
		wait for Clk_period;
		Addr <=  "00010000101010";
		Trees_din <= x"006710b1";
		wait for Clk_period;
		Addr <=  "00010000101011";
		Trees_din <= x"ff9210b1";
		wait for Clk_period;
		Addr <=  "00010000101100";
		Trees_din <= x"03fb1e0c";
		wait for Clk_period;
		Addr <=  "00010000101101";
		Trees_din <= x"0215a808";
		wait for Clk_period;
		Addr <=  "00010000101110";
		Trees_din <= x"00ff7304";
		wait for Clk_period;
		Addr <=  "00010000101111";
		Trees_din <= x"fff5112d";
		wait for Clk_period;
		Addr <=  "00010000110000";
		Trees_din <= x"ff6a112d";
		wait for Clk_period;
		Addr <=  "00010000110001";
		Trees_din <= x"003b112d";
		wait for Clk_period;
		Addr <=  "00010000110010";
		Trees_din <= x"04fd5308";
		wait for Clk_period;
		Addr <=  "00010000110011";
		Trees_din <= x"1b004804";
		wait for Clk_period;
		Addr <=  "00010000110100";
		Trees_din <= x"ff77112d";
		wait for Clk_period;
		Addr <=  "00010000110101";
		Trees_din <= x"0045112d";
		wait for Clk_period;
		Addr <=  "00010000110110";
		Trees_din <= x"040e641c";
		wait for Clk_period;
		Addr <=  "00010000110111";
		Trees_din <= x"1600010c";
		wait for Clk_period;
		Addr <=  "00010000111000";
		Trees_din <= x"15009504";
		wait for Clk_period;
		Addr <=  "00010000111001";
		Trees_din <= x"ffcf112d";
		wait for Clk_period;
		Addr <=  "00010000111010";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00010000111011";
		Trees_din <= x"00ae112d";
		wait for Clk_period;
		Addr <=  "00010000111100";
		Trees_din <= x"0038112d";
		wait for Clk_period;
		Addr <=  "00010000111101";
		Trees_din <= x"07005a08";
		wait for Clk_period;
		Addr <=  "00010000111110";
		Trees_din <= x"0c03e204";
		wait for Clk_period;
		Addr <=  "00010000111111";
		Trees_din <= x"0001112d";
		wait for Clk_period;
		Addr <=  "00010001000000";
		Trees_din <= x"007d112d";
		wait for Clk_period;
		Addr <=  "00010001000001";
		Trees_din <= x"0afa9a04";
		wait for Clk_period;
		Addr <=  "00010001000010";
		Trees_din <= x"0040112d";
		wait for Clk_period;
		Addr <=  "00010001000011";
		Trees_din <= x"ffb3112d";
		wait for Clk_period;
		Addr <=  "00010001000100";
		Trees_din <= x"05f9530c";
		wait for Clk_period;
		Addr <=  "00010001000101";
		Trees_din <= x"0f00b304";
		wait for Clk_period;
		Addr <=  "00010001000110";
		Trees_din <= x"006b112d";
		wait for Clk_period;
		Addr <=  "00010001000111";
		Trees_din <= x"0800ba04";
		wait for Clk_period;
		Addr <=  "00010001001000";
		Trees_din <= x"ff91112d";
		wait for Clk_period;
		Addr <=  "00010001001001";
		Trees_din <= x"0012112d";
		wait for Clk_period;
		Addr <=  "00010001001010";
		Trees_din <= x"008a112d";
		wait for Clk_period;
		Addr <=  "00010001001011";
		Trees_din <= x"03fb1e0c";
		wait for Clk_period;
		Addr <=  "00010001001100";
		Trees_din <= x"1c005008";
		wait for Clk_period;
		Addr <=  "00010001001101";
		Trees_din <= x"00ff7304";
		wait for Clk_period;
		Addr <=  "00010001001110";
		Trees_din <= x"fff111b9";
		wait for Clk_period;
		Addr <=  "00010001001111";
		Trees_din <= x"ff6b11b9";
		wait for Clk_period;
		Addr <=  "00010001010000";
		Trees_din <= x"004811b9";
		wait for Clk_period;
		Addr <=  "00010001010001";
		Trees_din <= x"04fd5308";
		wait for Clk_period;
		Addr <=  "00010001010010";
		Trees_din <= x"1500ae04";
		wait for Clk_period;
		Addr <=  "00010001010011";
		Trees_din <= x"ff7a11b9";
		wait for Clk_period;
		Addr <=  "00010001010100";
		Trees_din <= x"004111b9";
		wait for Clk_period;
		Addr <=  "00010001010101";
		Trees_din <= x"040a4a18";
		wait for Clk_period;
		Addr <=  "00010001010110";
		Trees_din <= x"1d003608";
		wait for Clk_period;
		Addr <=  "00010001010111";
		Trees_din <= x"11006c04";
		wait for Clk_period;
		Addr <=  "00010001011000";
		Trees_din <= x"001c11b9";
		wait for Clk_period;
		Addr <=  "00010001011001";
		Trees_din <= x"ff6711b9";
		wait for Clk_period;
		Addr <=  "00010001011010";
		Trees_din <= x"18003c08";
		wait for Clk_period;
		Addr <=  "00010001011011";
		Trees_din <= x"0c013804";
		wait for Clk_period;
		Addr <=  "00010001011100";
		Trees_din <= x"008611b9";
		wait for Clk_period;
		Addr <=  "00010001011101";
		Trees_din <= x"000011b9";
		wait for Clk_period;
		Addr <=  "00010001011110";
		Trees_din <= x"1d004204";
		wait for Clk_period;
		Addr <=  "00010001011111";
		Trees_din <= x"ffac11b9";
		wait for Clk_period;
		Addr <=  "00010001100000";
		Trees_din <= x"000211b9";
		wait for Clk_period;
		Addr <=  "00010001100001";
		Trees_din <= x"0700550c";
		wait for Clk_period;
		Addr <=  "00010001100010";
		Trees_din <= x"0bf98b04";
		wait for Clk_period;
		Addr <=  "00010001100011";
		Trees_din <= x"ffc611b9";
		wait for Clk_period;
		Addr <=  "00010001100100";
		Trees_din <= x"06f2a604";
		wait for Clk_period;
		Addr <=  "00010001100101";
		Trees_din <= x"002411b9";
		wait for Clk_period;
		Addr <=  "00010001100110";
		Trees_din <= x"00a811b9";
		wait for Clk_period;
		Addr <=  "00010001100111";
		Trees_din <= x"08000908";
		wait for Clk_period;
		Addr <=  "00010001101000";
		Trees_din <= x"09005604";
		wait for Clk_period;
		Addr <=  "00010001101001";
		Trees_din <= x"fffc11b9";
		wait for Clk_period;
		Addr <=  "00010001101010";
		Trees_din <= x"ff5c11b9";
		wait for Clk_period;
		Addr <=  "00010001101011";
		Trees_din <= x"0afccf04";
		wait for Clk_period;
		Addr <=  "00010001101100";
		Trees_din <= x"006611b9";
		wait for Clk_period;
		Addr <=  "00010001101101";
		Trees_din <= x"ffed11b9";
		wait for Clk_period;
		Addr <=  "00010001101110";
		Trees_din <= x"03fb1e0c";
		wait for Clk_period;
		Addr <=  "00010001101111";
		Trees_din <= x"1c005008";
		wait for Clk_period;
		Addr <=  "00010001110000";
		Trees_din <= x"00ff7304";
		wait for Clk_period;
		Addr <=  "00010001110001";
		Trees_din <= x"fff5124d";
		wait for Clk_period;
		Addr <=  "00010001110010";
		Trees_din <= x"ff6d124d";
		wait for Clk_period;
		Addr <=  "00010001110011";
		Trees_din <= x"0044124d";
		wait for Clk_period;
		Addr <=  "00010001110100";
		Trees_din <= x"06fa5b38";
		wait for Clk_period;
		Addr <=  "00010001110101";
		Trees_din <= x"0d039d20";
		wait for Clk_period;
		Addr <=  "00010001110110";
		Trees_din <= x"17000010";
		wait for Clk_period;
		Addr <=  "00010001110111";
		Trees_din <= x"16012208";
		wait for Clk_period;
		Addr <=  "00010001111000";
		Trees_din <= x"12fd8104";
		wait for Clk_period;
		Addr <=  "00010001111001";
		Trees_din <= x"ff93124d";
		wait for Clk_period;
		Addr <=  "00010001111010";
		Trees_din <= x"003a124d";
		wait for Clk_period;
		Addr <=  "00010001111011";
		Trees_din <= x"04086a04";
		wait for Clk_period;
		Addr <=  "00010001111100";
		Trees_din <= x"ff70124d";
		wait for Clk_period;
		Addr <=  "00010001111101";
		Trees_din <= x"0041124d";
		wait for Clk_period;
		Addr <=  "00010001111110";
		Trees_din <= x"14036408";
		wait for Clk_period;
		Addr <=  "00010001111111";
		Trees_din <= x"1c002504";
		wait for Clk_period;
		Addr <=  "00010010000000";
		Trees_din <= x"ffa3124d";
		wait for Clk_period;
		Addr <=  "00010010000001";
		Trees_din <= x"0003124d";
		wait for Clk_period;
		Addr <=  "00010010000010";
		Trees_din <= x"05fdfd04";
		wait for Clk_period;
		Addr <=  "00010010000011";
		Trees_din <= x"ff5e124d";
		wait for Clk_period;
		Addr <=  "00010010000100";
		Trees_din <= x"fffd124d";
		wait for Clk_period;
		Addr <=  "00010010000101";
		Trees_din <= x"0900550c";
		wait for Clk_period;
		Addr <=  "00010010000110";
		Trees_din <= x"13ffc108";
		wait for Clk_period;
		Addr <=  "00010010000111";
		Trees_din <= x"12fffc04";
		wait for Clk_period;
		Addr <=  "00010010001000";
		Trees_din <= x"fff1124d";
		wait for Clk_period;
		Addr <=  "00010010001001";
		Trees_din <= x"00a3124d";
		wait for Clk_period;
		Addr <=  "00010010001010";
		Trees_din <= x"ffdb124d";
		wait for Clk_period;
		Addr <=  "00010010001011";
		Trees_din <= x"0e03b208";
		wait for Clk_period;
		Addr <=  "00010010001100";
		Trees_din <= x"040c1204";
		wait for Clk_period;
		Addr <=  "00010010001101";
		Trees_din <= x"ff7b124d";
		wait for Clk_period;
		Addr <=  "00010010001110";
		Trees_din <= x"003c124d";
		wait for Clk_period;
		Addr <=  "00010010001111";
		Trees_din <= x"0077124d";
		wait for Clk_period;
		Addr <=  "00010010010000";
		Trees_din <= x"0c033d04";
		wait for Clk_period;
		Addr <=  "00010010010001";
		Trees_din <= x"ff81124d";
		wait for Clk_period;
		Addr <=  "00010010010010";
		Trees_din <= x"ffea124d";
		wait for Clk_period;
		Addr <=  "00010010010011";
		Trees_din <= x"00097444";
		wait for Clk_period;
		Addr <=  "00010010010100";
		Trees_din <= x"040c1228";
		wait for Clk_period;
		Addr <=  "00010010010101";
		Trees_din <= x"1d003508";
		wait for Clk_period;
		Addr <=  "00010010010110";
		Trees_din <= x"11006c04";
		wait for Clk_period;
		Addr <=  "00010010010111";
		Trees_din <= x"001812e9";
		wait for Clk_period;
		Addr <=  "00010010011000";
		Trees_din <= x"ff7012e9";
		wait for Clk_period;
		Addr <=  "00010010011001";
		Trees_din <= x"05fcb210";
		wait for Clk_period;
		Addr <=  "00010010011010";
		Trees_din <= x"05fc6908";
		wait for Clk_period;
		Addr <=  "00010010011011";
		Trees_din <= x"00037704";
		wait for Clk_period;
		Addr <=  "00010010011100";
		Trees_din <= x"000912e9";
		wait for Clk_period;
		Addr <=  "00010010011101";
		Trees_din <= x"ff9312e9";
		wait for Clk_period;
		Addr <=  "00010010011110";
		Trees_din <= x"0c00cd04";
		wait for Clk_period;
		Addr <=  "00010010011111";
		Trees_din <= x"000212e9";
		wait for Clk_period;
		Addr <=  "00010010100000";
		Trees_din <= x"ff3e12e9";
		wait for Clk_period;
		Addr <=  "00010010100001";
		Trees_din <= x"1d005608";
		wait for Clk_period;
		Addr <=  "00010010100010";
		Trees_din <= x"1a00b904";
		wait for Clk_period;
		Addr <=  "00010010100011";
		Trees_din <= x"ffb912e9";
		wait for Clk_period;
		Addr <=  "00010010100100";
		Trees_din <= x"002912e9";
		wait for Clk_period;
		Addr <=  "00010010100101";
		Trees_din <= x"1e009304";
		wait for Clk_period;
		Addr <=  "00010010100110";
		Trees_din <= x"00ec12e9";
		wait for Clk_period;
		Addr <=  "00010010100111";
		Trees_din <= x"001512e9";
		wait for Clk_period;
		Addr <=  "00010010101000";
		Trees_din <= x"07005504";
		wait for Clk_period;
		Addr <=  "00010010101001";
		Trees_din <= x"008412e9";
		wait for Clk_period;
		Addr <=  "00010010101010";
		Trees_din <= x"12fe6c08";
		wait for Clk_period;
		Addr <=  "00010010101011";
		Trees_din <= x"05fac804";
		wait for Clk_period;
		Addr <=  "00010010101100";
		Trees_din <= x"ff7912e9";
		wait for Clk_period;
		Addr <=  "00010010101101";
		Trees_din <= x"ffeb12e9";
		wait for Clk_period;
		Addr <=  "00010010101110";
		Trees_din <= x"05f89408";
		wait for Clk_period;
		Addr <=  "00010010101111";
		Trees_din <= x"0200af04";
		wait for Clk_period;
		Addr <=  "00010010110000";
		Trees_din <= x"000812e9";
		wait for Clk_period;
		Addr <=  "00010010110001";
		Trees_din <= x"ff9712e9";
		wait for Clk_period;
		Addr <=  "00010010110010";
		Trees_din <= x"02fac504";
		wait for Clk_period;
		Addr <=  "00010010110011";
		Trees_din <= x"ffb812e9";
		wait for Clk_period;
		Addr <=  "00010010110100";
		Trees_din <= x"007a12e9";
		wait for Clk_period;
		Addr <=  "00010010110101";
		Trees_din <= x"0e04b108";
		wait for Clk_period;
		Addr <=  "00010010110110";
		Trees_din <= x"05f70004";
		wait for Clk_period;
		Addr <=  "00010010110111";
		Trees_din <= x"003512e9";
		wait for Clk_period;
		Addr <=  "00010010111000";
		Trees_din <= x"ff6e12e9";
		wait for Clk_period;
		Addr <=  "00010010111001";
		Trees_din <= x"002412e9";
		wait for Clk_period;
		Addr <=  "00010010111010";
		Trees_din <= x"04faa904";
		wait for Clk_period;
		Addr <=  "00010010111011";
		Trees_din <= x"ff72136d";
		wait for Clk_period;
		Addr <=  "00010010111100";
		Trees_din <= x"03fb1e0c";
		wait for Clk_period;
		Addr <=  "00010010111101";
		Trees_din <= x"1d005408";
		wait for Clk_period;
		Addr <=  "00010010111110";
		Trees_din <= x"00ff7304";
		wait for Clk_period;
		Addr <=  "00010010111111";
		Trees_din <= x"ffda136d";
		wait for Clk_period;
		Addr <=  "00010011000000";
		Trees_din <= x"ff7b136d";
		wait for Clk_period;
		Addr <=  "00010011000001";
		Trees_din <= x"006c136d";
		wait for Clk_period;
		Addr <=  "00010011000010";
		Trees_din <= x"0d039d1c";
		wait for Clk_period;
		Addr <=  "00010011000011";
		Trees_din <= x"0c00610c";
		wait for Clk_period;
		Addr <=  "00010011000100";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00010011000101";
		Trees_din <= x"ff91136d";
		wait for Clk_period;
		Addr <=  "00010011000110";
		Trees_din <= x"1f000004";
		wait for Clk_period;
		Addr <=  "00010011000111";
		Trees_din <= x"0067136d";
		wait for Clk_period;
		Addr <=  "00010011001000";
		Trees_din <= x"ff92136d";
		wait for Clk_period;
		Addr <=  "00010011001001";
		Trees_din <= x"07005608";
		wait for Clk_period;
		Addr <=  "00010011001010";
		Trees_din <= x"06f7f304";
		wait for Clk_period;
		Addr <=  "00010011001011";
		Trees_din <= x"001d136d";
		wait for Clk_period;
		Addr <=  "00010011001100";
		Trees_din <= x"ff93136d";
		wait for Clk_period;
		Addr <=  "00010011001101";
		Trees_din <= x"1104ca04";
		wait for Clk_period;
		Addr <=  "00010011001110";
		Trees_din <= x"ffd3136d";
		wait for Clk_period;
		Addr <=  "00010011001111";
		Trees_din <= x"006f136d";
		wait for Clk_period;
		Addr <=  "00010011010000";
		Trees_din <= x"0900530c";
		wait for Clk_period;
		Addr <=  "00010011010001";
		Trees_din <= x"18004b08";
		wait for Clk_period;
		Addr <=  "00010011010010";
		Trees_din <= x"0f003204";
		wait for Clk_period;
		Addr <=  "00010011010011";
		Trees_din <= x"002a136d";
		wait for Clk_period;
		Addr <=  "00010011010100";
		Trees_din <= x"00b2136d";
		wait for Clk_period;
		Addr <=  "00010011010101";
		Trees_din <= x"ffc9136d";
		wait for Clk_period;
		Addr <=  "00010011010110";
		Trees_din <= x"0e03b208";
		wait for Clk_period;
		Addr <=  "00010011010111";
		Trees_din <= x"04086a04";
		wait for Clk_period;
		Addr <=  "00010011011000";
		Trees_din <= x"ff80136d";
		wait for Clk_period;
		Addr <=  "00010011011001";
		Trees_din <= x"0027136d";
		wait for Clk_period;
		Addr <=  "00010011011010";
		Trees_din <= x"0076136d";
		wait for Clk_period;
		Addr <=  "00010011011011";
		Trees_din <= x"04faa904";
		wait for Clk_period;
		Addr <=  "00010011011100";
		Trees_din <= x"ff7413e1";
		wait for Clk_period;
		Addr <=  "00010011011101";
		Trees_din <= x"040e642c";
		wait for Clk_period;
		Addr <=  "00010011011110";
		Trees_din <= x"0afb0b14";
		wait for Clk_period;
		Addr <=  "00010011011111";
		Trees_din <= x"0eff2d04";
		wait for Clk_period;
		Addr <=  "00010011100000";
		Trees_din <= x"010213e1";
		wait for Clk_period;
		Addr <=  "00010011100001";
		Trees_din <= x"0301f908";
		wait for Clk_period;
		Addr <=  "00010011100010";
		Trees_din <= x"15008d04";
		wait for Clk_period;
		Addr <=  "00010011100011";
		Trees_din <= x"004e13e1";
		wait for Clk_period;
		Addr <=  "00010011100100";
		Trees_din <= x"ff9513e1";
		wait for Clk_period;
		Addr <=  "00010011100101";
		Trees_din <= x"06f7dd04";
		wait for Clk_period;
		Addr <=  "00010011100110";
		Trees_din <= x"006313e1";
		wait for Clk_period;
		Addr <=  "00010011100111";
		Trees_din <= x"ffc613e1";
		wait for Clk_period;
		Addr <=  "00010011101000";
		Trees_din <= x"04fff308";
		wait for Clk_period;
		Addr <=  "00010011101001";
		Trees_din <= x"0e04b104";
		wait for Clk_period;
		Addr <=  "00010011101010";
		Trees_din <= x"ff7613e1";
		wait for Clk_period;
		Addr <=  "00010011101011";
		Trees_din <= x"003a13e1";
		wait for Clk_period;
		Addr <=  "00010011101100";
		Trees_din <= x"05fcb208";
		wait for Clk_period;
		Addr <=  "00010011101101";
		Trees_din <= x"05fc1204";
		wait for Clk_period;
		Addr <=  "00010011101110";
		Trees_din <= x"fff713e1";
		wait for Clk_period;
		Addr <=  "00010011101111";
		Trees_din <= x"ff8d13e1";
		wait for Clk_period;
		Addr <=  "00010011110000";
		Trees_din <= x"1700de04";
		wait for Clk_period;
		Addr <=  "00010011110001";
		Trees_din <= x"003013e1";
		wait for Clk_period;
		Addr <=  "00010011110010";
		Trees_din <= x"ffd713e1";
		wait for Clk_period;
		Addr <=  "00010011110011";
		Trees_din <= x"09005408";
		wait for Clk_period;
		Addr <=  "00010011110100";
		Trees_din <= x"06f16a04";
		wait for Clk_period;
		Addr <=  "00010011110101";
		Trees_din <= x"ffce13e1";
		wait for Clk_period;
		Addr <=  "00010011110110";
		Trees_din <= x"005913e1";
		wait for Clk_period;
		Addr <=  "00010011110111";
		Trees_din <= x"007813e1";
		wait for Clk_period;
		Addr <=  "00010011111000";
		Trees_din <= x"04faa904";
		wait for Clk_period;
		Addr <=  "00010011111001";
		Trees_din <= x"ff771455";
		wait for Clk_period;
		Addr <=  "00010011111010";
		Trees_din <= x"010de930";
		wait for Clk_period;
		Addr <=  "00010011111011";
		Trees_din <= x"1a008e10";
		wait for Clk_period;
		Addr <=  "00010011111100";
		Trees_din <= x"0bfa9f04";
		wait for Clk_period;
		Addr <=  "00010011111101";
		Trees_din <= x"ffa01455";
		wait for Clk_period;
		Addr <=  "00010011111110";
		Trees_din <= x"08009d08";
		wait for Clk_period;
		Addr <=  "00010011111111";
		Trees_din <= x"01fc5904";
		wait for Clk_period;
		Addr <=  "00010100000000";
		Trees_din <= x"00681455";
		wait for Clk_period;
		Addr <=  "00010100000001";
		Trees_din <= x"ffd51455";
		wait for Clk_period;
		Addr <=  "00010100000010";
		Trees_din <= x"00d11455";
		wait for Clk_period;
		Addr <=  "00010100000011";
		Trees_din <= x"040a4a10";
		wait for Clk_period;
		Addr <=  "00010100000100";
		Trees_din <= x"18004b08";
		wait for Clk_period;
		Addr <=  "00010100000101";
		Trees_din <= x"0f006404";
		wait for Clk_period;
		Addr <=  "00010100000110";
		Trees_din <= x"00221455";
		wait for Clk_period;
		Addr <=  "00010100000111";
		Trees_din <= x"ffe81455";
		wait for Clk_period;
		Addr <=  "00010100001000";
		Trees_din <= x"0bfad604";
		wait for Clk_period;
		Addr <=  "00010100001001";
		Trees_din <= x"00361455";
		wait for Clk_period;
		Addr <=  "00010100001010";
		Trees_din <= x"ff711455";
		wait for Clk_period;
		Addr <=  "00010100001011";
		Trees_din <= x"07005508";
		wait for Clk_period;
		Addr <=  "00010100001100";
		Trees_din <= x"0bf98b04";
		wait for Clk_period;
		Addr <=  "00010100001101";
		Trees_din <= x"ffca1455";
		wait for Clk_period;
		Addr <=  "00010100001110";
		Trees_din <= x"007a1455";
		wait for Clk_period;
		Addr <=  "00010100001111";
		Trees_din <= x"12fe6c04";
		wait for Clk_period;
		Addr <=  "00010100010000";
		Trees_din <= x"ffa91455";
		wait for Clk_period;
		Addr <=  "00010100010001";
		Trees_din <= x"00181455";
		wait for Clk_period;
		Addr <=  "00010100010010";
		Trees_din <= x"0b048204";
		wait for Clk_period;
		Addr <=  "00010100010011";
		Trees_din <= x"ff841455";
		wait for Clk_period;
		Addr <=  "00010100010100";
		Trees_din <= x"00141455";
		wait for Clk_period;
		Addr <=  "00010100010101";
		Trees_din <= x"03fb1e0c";
		wait for Clk_period;
		Addr <=  "00010100010110";
		Trees_din <= x"1d005408";
		wait for Clk_period;
		Addr <=  "00010100010111";
		Trees_din <= x"1900ac04";
		wait for Clk_period;
		Addr <=  "00010100011000";
		Trees_din <= x"ff7514d1";
		wait for Clk_period;
		Addr <=  "00010100011001";
		Trees_din <= x"ffd914d1";
		wait for Clk_period;
		Addr <=  "00010100011010";
		Trees_din <= x"002514d1";
		wait for Clk_period;
		Addr <=  "00010100011011";
		Trees_din <= x"0d039d18";
		wait for Clk_period;
		Addr <=  "00010100011100";
		Trees_din <= x"04fd5304";
		wait for Clk_period;
		Addr <=  "00010100011101";
		Trees_din <= x"ff8914d1";
		wait for Clk_period;
		Addr <=  "00010100011110";
		Trees_din <= x"10f72e04";
		wait for Clk_period;
		Addr <=  "00010100011111";
		Trees_din <= x"ff7e14d1";
		wait for Clk_period;
		Addr <=  "00010100100000";
		Trees_din <= x"05f8b408";
		wait for Clk_period;
		Addr <=  "00010100100001";
		Trees_din <= x"11fdfc04";
		wait for Clk_period;
		Addr <=  "00010100100010";
		Trees_din <= x"005714d1";
		wait for Clk_period;
		Addr <=  "00010100100011";
		Trees_din <= x"ff9f14d1";
		wait for Clk_period;
		Addr <=  "00010100100100";
		Trees_din <= x"1c002504";
		wait for Clk_period;
		Addr <=  "00010100100101";
		Trees_din <= x"ffad14d1";
		wait for Clk_period;
		Addr <=  "00010100100110";
		Trees_din <= x"000e14d1";
		wait for Clk_period;
		Addr <=  "00010100100111";
		Trees_din <= x"09005310";
		wait for Clk_period;
		Addr <=  "00010100101000";
		Trees_din <= x"1102f10c";
		wait for Clk_period;
		Addr <=  "00010100101001";
		Trees_din <= x"1b004908";
		wait for Clk_period;
		Addr <=  "00010100101010";
		Trees_din <= x"0b048504";
		wait for Clk_period;
		Addr <=  "00010100101011";
		Trees_din <= x"00ae14d1";
		wait for Clk_period;
		Addr <=  "00010100101100";
		Trees_din <= x"003b14d1";
		wait for Clk_period;
		Addr <=  "00010100101101";
		Trees_din <= x"ffe814d1";
		wait for Clk_period;
		Addr <=  "00010100101110";
		Trees_din <= x"ffc614d1";
		wait for Clk_period;
		Addr <=  "00010100101111";
		Trees_din <= x"0e03b508";
		wait for Clk_period;
		Addr <=  "00010100110000";
		Trees_din <= x"0409d604";
		wait for Clk_period;
		Addr <=  "00010100110001";
		Trees_din <= x"ff8614d1";
		wait for Clk_period;
		Addr <=  "00010100110010";
		Trees_din <= x"002314d1";
		wait for Clk_period;
		Addr <=  "00010100110011";
		Trees_din <= x"006514d1";
		wait for Clk_period;
		Addr <=  "00010100110100";
		Trees_din <= x"04faa904";
		wait for Clk_period;
		Addr <=  "00010100110101";
		Trees_din <= x"ff7c1515";
		wait for Clk_period;
		Addr <=  "00010100110110";
		Trees_din <= x"04fac204";
		wait for Clk_period;
		Addr <=  "00010100110111";
		Trees_din <= x"00b81515";
		wait for Clk_period;
		Addr <=  "00010100111000";
		Trees_din <= x"03fb1e08";
		wait for Clk_period;
		Addr <=  "00010100111001";
		Trees_din <= x"00ff7304";
		wait for Clk_period;
		Addr <=  "00010100111010";
		Trees_din <= x"fffa1515";
		wait for Clk_period;
		Addr <=  "00010100111011";
		Trees_din <= x"ff831515";
		wait for Clk_period;
		Addr <=  "00010100111100";
		Trees_din <= x"0ef8ef04";
		wait for Clk_period;
		Addr <=  "00010100111101";
		Trees_din <= x"ff921515";
		wait for Clk_period;
		Addr <=  "00010100111110";
		Trees_din <= x"040e6408";
		wait for Clk_period;
		Addr <=  "00010100111111";
		Trees_din <= x"0efe0804";
		wait for Clk_period;
		Addr <=  "00010101000000";
		Trees_din <= x"00211515";
		wait for Clk_period;
		Addr <=  "00010101000001";
		Trees_din <= x"fff71515";
		wait for Clk_period;
		Addr <=  "00010101000010";
		Trees_din <= x"00fd6404";
		wait for Clk_period;
		Addr <=  "00010101000011";
		Trees_din <= x"006b1515";
		wait for Clk_period;
		Addr <=  "00010101000100";
		Trees_din <= x"fffc1515";
		wait for Clk_period;
		Addr <=  "00010101000101";
		Trees_din <= x"04faa904";
		wait for Clk_period;
		Addr <=  "00010101000110";
		Trees_din <= x"ff7f1561";
		wait for Clk_period;
		Addr <=  "00010101000111";
		Trees_din <= x"04fac204";
		wait for Clk_period;
		Addr <=  "00010101001000";
		Trees_din <= x"00a61561";
		wait for Clk_period;
		Addr <=  "00010101001001";
		Trees_din <= x"04fd5304";
		wait for Clk_period;
		Addr <=  "00010101001010";
		Trees_din <= x"ff891561";
		wait for Clk_period;
		Addr <=  "00010101001011";
		Trees_din <= x"040e6410";
		wait for Clk_period;
		Addr <=  "00010101001100";
		Trees_din <= x"06f44e08";
		wait for Clk_period;
		Addr <=  "00010101001101";
		Trees_din <= x"0afccf04";
		wait for Clk_period;
		Addr <=  "00010101001110";
		Trees_din <= x"000d1561";
		wait for Clk_period;
		Addr <=  "00010101001111";
		Trees_din <= x"ffbc1561";
		wait for Clk_period;
		Addr <=  "00010101010000";
		Trees_din <= x"1a00fe04";
		wait for Clk_period;
		Addr <=  "00010101010001";
		Trees_din <= x"00101561";
		wait for Clk_period;
		Addr <=  "00010101010010";
		Trees_din <= x"ffa51561";
		wait for Clk_period;
		Addr <=  "00010101010011";
		Trees_din <= x"05f95308";
		wait for Clk_period;
		Addr <=  "00010101010100";
		Trees_din <= x"0f00b304";
		wait for Clk_period;
		Addr <=  "00010101010101";
		Trees_din <= x"00511561";
		wait for Clk_period;
		Addr <=  "00010101010110";
		Trees_din <= x"ffc71561";
		wait for Clk_period;
		Addr <=  "00010101010111";
		Trees_din <= x"00761561";
		wait for Clk_period;
		Addr <=  "00010101011000";
		Trees_din <= x"00097438";
		wait for Clk_period;
		Addr <=  "00010101011001";
		Trees_din <= x"10058f28";
		wait for Clk_period;
		Addr <=  "00010101011010";
		Trees_din <= x"1005591c";
		wait for Clk_period;
		Addr <=  "00010101011011";
		Trees_din <= x"1a008e0c";
		wait for Clk_period;
		Addr <=  "00010101011100";
		Trees_din <= x"0e00b808";
		wait for Clk_period;
		Addr <=  "00010101011101";
		Trees_din <= x"1200e704";
		wait for Clk_period;
		Addr <=  "00010101011110";
		Trees_din <= x"002715e5";
		wait for Clk_period;
		Addr <=  "00010101011111";
		Trees_din <= x"00ad15e5";
		wait for Clk_period;
		Addr <=  "00010101100000";
		Trees_din <= x"ffeb15e5";
		wait for Clk_period;
		Addr <=  "00010101100001";
		Trees_din <= x"1200c308";
		wait for Clk_period;
		Addr <=  "00010101100010";
		Trees_din <= x"12fda004";
		wait for Clk_period;
		Addr <=  "00010101100011";
		Trees_din <= x"ffce15e5";
		wait for Clk_period;
		Addr <=  "00010101100100";
		Trees_din <= x"002d15e5";
		wait for Clk_period;
		Addr <=  "00010101100101";
		Trees_din <= x"10f95704";
		wait for Clk_period;
		Addr <=  "00010101100110";
		Trees_din <= x"ff9915e5";
		wait for Clk_period;
		Addr <=  "00010101100111";
		Trees_din <= x"fff815e5";
		wait for Clk_period;
		Addr <=  "00010101101000";
		Trees_din <= x"0afb2e04";
		wait for Clk_period;
		Addr <=  "00010101101001";
		Trees_din <= x"008815e5";
		wait for Clk_period;
		Addr <=  "00010101101010";
		Trees_din <= x"07005804";
		wait for Clk_period;
		Addr <=  "00010101101011";
		Trees_din <= x"ffa915e5";
		wait for Clk_period;
		Addr <=  "00010101101100";
		Trees_din <= x"003f15e5";
		wait for Clk_period;
		Addr <=  "00010101101101";
		Trees_din <= x"0d01d90c";
		wait for Clk_period;
		Addr <=  "00010101101110";
		Trees_din <= x"01030e08";
		wait for Clk_period;
		Addr <=  "00010101101111";
		Trees_din <= x"09005704";
		wait for Clk_period;
		Addr <=  "00010101110000";
		Trees_din <= x"006f15e5";
		wait for Clk_period;
		Addr <=  "00010101110001";
		Trees_din <= x"ffe515e5";
		wait for Clk_period;
		Addr <=  "00010101110010";
		Trees_din <= x"ff9a15e5";
		wait for Clk_period;
		Addr <=  "00010101110011";
		Trees_din <= x"ff8115e5";
		wait for Clk_period;
		Addr <=  "00010101110100";
		Trees_din <= x"1d003d08";
		wait for Clk_period;
		Addr <=  "00010101110101";
		Trees_din <= x"1900a404";
		wait for Clk_period;
		Addr <=  "00010101110110";
		Trees_din <= x"005d15e5";
		wait for Clk_period;
		Addr <=  "00010101110111";
		Trees_din <= x"ffa415e5";
		wait for Clk_period;
		Addr <=  "00010101111000";
		Trees_din <= x"ff7a15e5";
		wait for Clk_period;
		Addr <=  "00010101111001";
		Trees_din <= x"04faa904";
		wait for Clk_period;
		Addr <=  "00010101111010";
		Trees_din <= x"ff851629";
		wait for Clk_period;
		Addr <=  "00010101111011";
		Trees_din <= x"04fac204";
		wait for Clk_period;
		Addr <=  "00010101111100";
		Trees_din <= x"008c1629";
		wait for Clk_period;
		Addr <=  "00010101111101";
		Trees_din <= x"03fb1e08";
		wait for Clk_period;
		Addr <=  "00010101111110";
		Trees_din <= x"00ff7304";
		wait for Clk_period;
		Addr <=  "00010101111111";
		Trees_din <= x"fff71629";
		wait for Clk_period;
		Addr <=  "00010110000000";
		Trees_din <= x"ff8a1629";
		wait for Clk_period;
		Addr <=  "00010110000001";
		Trees_din <= x"0ef8ef04";
		wait for Clk_period;
		Addr <=  "00010110000010";
		Trees_din <= x"ff9e1629";
		wait for Clk_period;
		Addr <=  "00010110000011";
		Trees_din <= x"0404aa08";
		wait for Clk_period;
		Addr <=  "00010110000100";
		Trees_din <= x"06f4f204";
		wait for Clk_period;
		Addr <=  "00010110000101";
		Trees_din <= x"ff821629";
		wait for Clk_period;
		Addr <=  "00010110000110";
		Trees_din <= x"fffe1629";
		wait for Clk_period;
		Addr <=  "00010110000111";
		Trees_din <= x"0d034d04";
		wait for Clk_period;
		Addr <=  "00010110001000";
		Trees_din <= x"00031629";
		wait for Clk_period;
		Addr <=  "00010110001001";
		Trees_din <= x"003e1629";
		wait for Clk_period;
		Addr <=  "00010110001010";
		Trees_din <= x"04faa904";
		wait for Clk_period;
		Addr <=  "00010110001011";
		Trees_din <= x"ff881675";
		wait for Clk_period;
		Addr <=  "00010110001100";
		Trees_din <= x"04fac204";
		wait for Clk_period;
		Addr <=  "00010110001101";
		Trees_din <= x"007e1675";
		wait for Clk_period;
		Addr <=  "00010110001110";
		Trees_din <= x"04fd5304";
		wait for Clk_period;
		Addr <=  "00010110001111";
		Trees_din <= x"ff911675";
		wait for Clk_period;
		Addr <=  "00010110010000";
		Trees_din <= x"040c1210";
		wait for Clk_period;
		Addr <=  "00010110010001";
		Trees_din <= x"1d003508";
		wait for Clk_period;
		Addr <=  "00010110010010";
		Trees_din <= x"11015604";
		wait for Clk_period;
		Addr <=  "00010110010011";
		Trees_din <= x"fffe1675";
		wait for Clk_period;
		Addr <=  "00010110010100";
		Trees_din <= x"ff831675";
		wait for Clk_period;
		Addr <=  "00010110010101";
		Trees_din <= x"18003c04";
		wait for Clk_period;
		Addr <=  "00010110010110";
		Trees_din <= x"00231675";
		wait for Clk_period;
		Addr <=  "00010110010111";
		Trees_din <= x"fff11675";
		wait for Clk_period;
		Addr <=  "00010110011000";
		Trees_din <= x"07005504";
		wait for Clk_period;
		Addr <=  "00010110011001";
		Trees_din <= x"006e1675";
		wait for Clk_period;
		Addr <=  "00010110011010";
		Trees_din <= x"12fe6c04";
		wait for Clk_period;
		Addr <=  "00010110011011";
		Trees_din <= x"ffa71675";
		wait for Clk_period;
		Addr <=  "00010110011100";
		Trees_din <= x"002c1675";
		wait for Clk_period;
		Addr <=  "00010110011101";
		Trees_din <= x"04faa904";
		wait for Clk_period;
		Addr <=  "00010110011110";
		Trees_din <= x"ff8c16d1";
		wait for Clk_period;
		Addr <=  "00010110011111";
		Trees_din <= x"04fac204";
		wait for Clk_period;
		Addr <=  "00010110100000";
		Trees_din <= x"007416d1";
		wait for Clk_period;
		Addr <=  "00010110100001";
		Trees_din <= x"03fb1e08";
		wait for Clk_period;
		Addr <=  "00010110100010";
		Trees_din <= x"00011804";
		wait for Clk_period;
		Addr <=  "00010110100011";
		Trees_din <= x"fff116d1";
		wait for Clk_period;
		Addr <=  "00010110100100";
		Trees_din <= x"ff9016d1";
		wait for Clk_period;
		Addr <=  "00010110100101";
		Trees_din <= x"0206e310";
		wait for Clk_period;
		Addr <=  "00010110100110";
		Trees_din <= x"02055108";
		wait for Clk_period;
		Addr <=  "00010110100111";
		Trees_din <= x"0c004604";
		wait for Clk_period;
		Addr <=  "00010110101000";
		Trees_din <= x"003f16d1";
		wait for Clk_period;
		Addr <=  "00010110101001";
		Trees_din <= x"fffc16d1";
		wait for Clk_period;
		Addr <=  "00010110101010";
		Trees_din <= x"0802d604";
		wait for Clk_period;
		Addr <=  "00010110101011";
		Trees_din <= x"ff9616d1";
		wait for Clk_period;
		Addr <=  "00010110101100";
		Trees_din <= x"001f16d1";
		wait for Clk_period;
		Addr <=  "00010110101101";
		Trees_din <= x"0d025f08";
		wait for Clk_period;
		Addr <=  "00010110101110";
		Trees_din <= x"0d011004";
		wait for Clk_period;
		Addr <=  "00010110101111";
		Trees_din <= x"ffd016d1";
		wait for Clk_period;
		Addr <=  "00010110110000";
		Trees_din <= x"00b616d1";
		wait for Clk_period;
		Addr <=  "00010110110001";
		Trees_din <= x"08000c04";
		wait for Clk_period;
		Addr <=  "00010110110010";
		Trees_din <= x"003a16d1";
		wait for Clk_period;
		Addr <=  "00010110110011";
		Trees_din <= x"ff9516d1";
		wait for Clk_period;
		Addr <=  "00010110110100";
		Trees_din <= x"000c5848";
		wait for Clk_period;
		Addr <=  "00010110110101";
		Trees_din <= x"10058f38";
		wait for Clk_period;
		Addr <=  "00010110110110";
		Trees_din <= x"10050c20";
		wait for Clk_period;
		Addr <=  "00010110110111";
		Trees_din <= x"09005710";
		wait for Clk_period;
		Addr <=  "00010110111000";
		Trees_din <= x"06f42b08";
		wait for Clk_period;
		Addr <=  "00010110111001";
		Trees_din <= x"06f05e04";
		wait for Clk_period;
		Addr <=  "00010110111010";
		Trees_din <= x"0057176d";
		wait for Clk_period;
		Addr <=  "00010110111011";
		Trees_din <= x"ffca176d";
		wait for Clk_period;
		Addr <=  "00010110111100";
		Trees_din <= x"1a00f404";
		wait for Clk_period;
		Addr <=  "00010110111101";
		Trees_din <= x"002c176d";
		wait for Clk_period;
		Addr <=  "00010110111110";
		Trees_din <= x"ffc0176d";
		wait for Clk_period;
		Addr <=  "00010110111111";
		Trees_din <= x"06f37108";
		wait for Clk_period;
		Addr <=  "00010111000000";
		Trees_din <= x"15009704";
		wait for Clk_period;
		Addr <=  "00010111000001";
		Trees_din <= x"006d176d";
		wait for Clk_period;
		Addr <=  "00010111000010";
		Trees_din <= x"ffcd176d";
		wait for Clk_period;
		Addr <=  "00010111000011";
		Trees_din <= x"0a021e04";
		wait for Clk_period;
		Addr <=  "00010111000100";
		Trees_din <= x"ff8f176d";
		wait for Clk_period;
		Addr <=  "00010111000101";
		Trees_din <= x"fff1176d";
		wait for Clk_period;
		Addr <=  "00010111000110";
		Trees_din <= x"06f3bf08";
		wait for Clk_period;
		Addr <=  "00010111000111";
		Trees_din <= x"02013704";
		wait for Clk_period;
		Addr <=  "00010111001000";
		Trees_din <= x"0033176d";
		wait for Clk_period;
		Addr <=  "00010111001001";
		Trees_din <= x"ff7f176d";
		wait for Clk_period;
		Addr <=  "00010111001010";
		Trees_din <= x"04065f08";
		wait for Clk_period;
		Addr <=  "00010111001011";
		Trees_din <= x"02012d04";
		wait for Clk_period;
		Addr <=  "00010111001100";
		Trees_din <= x"ffba176d";
		wait for Clk_period;
		Addr <=  "00010111001101";
		Trees_din <= x"005a176d";
		wait for Clk_period;
		Addr <=  "00010111001110";
		Trees_din <= x"09004d04";
		wait for Clk_period;
		Addr <=  "00010111001111";
		Trees_din <= x"fff4176d";
		wait for Clk_period;
		Addr <=  "00010111010000";
		Trees_din <= x"00b0176d";
		wait for Clk_period;
		Addr <=  "00010111010001";
		Trees_din <= x"0d01d90c";
		wait for Clk_period;
		Addr <=  "00010111010010";
		Trees_din <= x"01030e08";
		wait for Clk_period;
		Addr <=  "00010111010011";
		Trees_din <= x"09005704";
		wait for Clk_period;
		Addr <=  "00010111010100";
		Trees_din <= x"005a176d";
		wait for Clk_period;
		Addr <=  "00010111010101";
		Trees_din <= x"ffe7176d";
		wait for Clk_period;
		Addr <=  "00010111010110";
		Trees_din <= x"ffa7176d";
		wait for Clk_period;
		Addr <=  "00010111010111";
		Trees_din <= x"ff8d176d";
		wait for Clk_period;
		Addr <=  "00010111011000";
		Trees_din <= x"05f8b404";
		wait for Clk_period;
		Addr <=  "00010111011001";
		Trees_din <= x"000e176d";
		wait for Clk_period;
		Addr <=  "00010111011010";
		Trees_din <= x"ff88176d";
		wait for Clk_period;
		Addr <=  "00010111011011";
		Trees_din <= x"0404aa34";
		wait for Clk_period;
		Addr <=  "00010111011100";
		Trees_din <= x"05fe701c";
		wait for Clk_period;
		Addr <=  "00010111011101";
		Trees_din <= x"1602f314";
		wait for Clk_period;
		Addr <=  "00010111011110";
		Trees_din <= x"0f005a08";
		wait for Clk_period;
		Addr <=  "00010111011111";
		Trees_din <= x"1a00d104";
		wait for Clk_period;
		Addr <=  "00010111100000";
		Trees_din <= x"ffca1861";
		wait for Clk_period;
		Addr <=  "00010111100001";
		Trees_din <= x"008a1861";
		wait for Clk_period;
		Addr <=  "00010111100010";
		Trees_din <= x"07005804";
		wait for Clk_period;
		Addr <=  "00010111100011";
		Trees_din <= x"ff7b1861";
		wait for Clk_period;
		Addr <=  "00010111100100";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00010111100101";
		Trees_din <= x"ffa41861";
		wait for Clk_period;
		Addr <=  "00010111100110";
		Trees_din <= x"004b1861";
		wait for Clk_period;
		Addr <=  "00010111100111";
		Trees_din <= x"05f8b404";
		wait for Clk_period;
		Addr <=  "00010111101000";
		Trees_din <= x"ffee1861";
		wait for Clk_period;
		Addr <=  "00010111101001";
		Trees_din <= x"ff761861";
		wait for Clk_period;
		Addr <=  "00010111101010";
		Trees_din <= x"0afb150c";
		wait for Clk_period;
		Addr <=  "00010111101011";
		Trees_din <= x"05fefa04";
		wait for Clk_period;
		Addr <=  "00010111101100";
		Trees_din <= x"00ab1861";
		wait for Clk_period;
		Addr <=  "00010111101101";
		Trees_din <= x"19008204";
		wait for Clk_period;
		Addr <=  "00010111101110";
		Trees_din <= x"006e1861";
		wait for Clk_period;
		Addr <=  "00010111101111";
		Trees_din <= x"ffc01861";
		wait for Clk_period;
		Addr <=  "00010111110000";
		Trees_din <= x"0efcb008";
		wait for Clk_period;
		Addr <=  "00010111110001";
		Trees_din <= x"0801fa04";
		wait for Clk_period;
		Addr <=  "00010111110010";
		Trees_din <= x"002a1861";
		wait for Clk_period;
		Addr <=  "00010111110011";
		Trees_din <= x"fff11861";
		wait for Clk_period;
		Addr <=  "00010111110100";
		Trees_din <= x"ffa01861";
		wait for Clk_period;
		Addr <=  "00010111110101";
		Trees_din <= x"0d034d2c";
		wait for Clk_period;
		Addr <=  "00010111110110";
		Trees_din <= x"0d02e11c";
		wait for Clk_period;
		Addr <=  "00010111110111";
		Trees_din <= x"08014810";
		wait for Clk_period;
		Addr <=  "00010111111000";
		Trees_din <= x"00fcaf08";
		wait for Clk_period;
		Addr <=  "00010111111001";
		Trees_din <= x"08000004";
		wait for Clk_period;
		Addr <=  "00010111111010";
		Trees_din <= x"ff931861";
		wait for Clk_period;
		Addr <=  "00010111111011";
		Trees_din <= x"003f1861";
		wait for Clk_period;
		Addr <=  "00010111111100";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00010111111101";
		Trees_din <= x"00361861";
		wait for Clk_period;
		Addr <=  "00010111111110";
		Trees_din <= x"ffaf1861";
		wait for Clk_period;
		Addr <=  "00010111111111";
		Trees_din <= x"07005b08";
		wait for Clk_period;
		Addr <=  "00011000000000";
		Trees_din <= x"01fe2604";
		wait for Clk_period;
		Addr <=  "00011000000001";
		Trees_din <= x"ffdd1861";
		wait for Clk_period;
		Addr <=  "00011000000010";
		Trees_din <= x"00571861";
		wait for Clk_period;
		Addr <=  "00011000000011";
		Trees_din <= x"ff981861";
		wait for Clk_period;
		Addr <=  "00011000000100";
		Trees_din <= x"1600f304";
		wait for Clk_period;
		Addr <=  "00011000000101";
		Trees_din <= x"00331861";
		wait for Clk_period;
		Addr <=  "00011000000110";
		Trees_din <= x"1500a808";
		wait for Clk_period;
		Addr <=  "00011000000111";
		Trees_din <= x"12003304";
		wait for Clk_period;
		Addr <=  "00011000001000";
		Trees_din <= x"ffdd1861";
		wait for Clk_period;
		Addr <=  "00011000001001";
		Trees_din <= x"ff621861";
		wait for Clk_period;
		Addr <=  "00011000001010";
		Trees_din <= x"001c1861";
		wait for Clk_period;
		Addr <=  "00011000001011";
		Trees_din <= x"0a02a214";
		wait for Clk_period;
		Addr <=  "00011000001100";
		Trees_din <= x"0409420c";
		wait for Clk_period;
		Addr <=  "00011000001101";
		Trees_din <= x"0f017f08";
		wait for Clk_period;
		Addr <=  "00011000001110";
		Trees_din <= x"09005504";
		wait for Clk_period;
		Addr <=  "00011000001111";
		Trees_din <= x"008a1861";
		wait for Clk_period;
		Addr <=  "00011000010000";
		Trees_din <= x"001b1861";
		wait for Clk_period;
		Addr <=  "00011000010001";
		Trees_din <= x"fff01861";
		wait for Clk_period;
		Addr <=  "00011000010010";
		Trees_din <= x"02fe4f04";
		wait for Clk_period;
		Addr <=  "00011000010011";
		Trees_din <= x"00281861";
		wait for Clk_period;
		Addr <=  "00011000010100";
		Trees_din <= x"ffce1861";
		wait for Clk_period;
		Addr <=  "00011000010101";
		Trees_din <= x"06f59704";
		wait for Clk_period;
		Addr <=  "00011000010110";
		Trees_din <= x"002e1861";
		wait for Clk_period;
		Addr <=  "00011000010111";
		Trees_din <= x"ffa71861";
		wait for Clk_period;
		Addr <=  "00011000011000";
		Trees_din <= x"000c5844";
		wait for Clk_period;
		Addr <=  "00011000011001";
		Trees_din <= x"040e643c";
		wait for Clk_period;
		Addr <=  "00011000011010";
		Trees_din <= x"06f41920";
		wait for Clk_period;
		Addr <=  "00011000011011";
		Trees_din <= x"0afccf10";
		wait for Clk_period;
		Addr <=  "00011000011100";
		Trees_din <= x"1101af08";
		wait for Clk_period;
		Addr <=  "00011000011101";
		Trees_din <= x"01071c04";
		wait for Clk_period;
		Addr <=  "00011000011110";
		Trees_din <= x"000818f5";
		wait for Clk_period;
		Addr <=  "00011000011111";
		Trees_din <= x"008918f5";
		wait for Clk_period;
		Addr <=  "00011000100000";
		Trees_din <= x"0afcba04";
		wait for Clk_period;
		Addr <=  "00011000100001";
		Trees_din <= x"ffaa18f5";
		wait for Clk_period;
		Addr <=  "00011000100010";
		Trees_din <= x"005318f5";
		wait for Clk_period;
		Addr <=  "00011000100011";
		Trees_din <= x"00fda608";
		wait for Clk_period;
		Addr <=  "00011000100100";
		Trees_din <= x"15009204";
		wait for Clk_period;
		Addr <=  "00011000100101";
		Trees_din <= x"ffad18f5";
		wait for Clk_period;
		Addr <=  "00011000100110";
		Trees_din <= x"003318f5";
		wait for Clk_period;
		Addr <=  "00011000100111";
		Trees_din <= x"02ff2a04";
		wait for Clk_period;
		Addr <=  "00011000101000";
		Trees_din <= x"fff518f5";
		wait for Clk_period;
		Addr <=  "00011000101001";
		Trees_din <= x"ff7718f5";
		wait for Clk_period;
		Addr <=  "00011000101010";
		Trees_din <= x"1d00380c";
		wait for Clk_period;
		Addr <=  "00011000101011";
		Trees_din <= x"0e03e108";
		wait for Clk_period;
		Addr <=  "00011000101100";
		Trees_din <= x"0afaf604";
		wait for Clk_period;
		Addr <=  "00011000101101";
		Trees_din <= x"000618f5";
		wait for Clk_period;
		Addr <=  "00011000101110";
		Trees_din <= x"ff7a18f5";
		wait for Clk_period;
		Addr <=  "00011000101111";
		Trees_din <= x"004b18f5";
		wait for Clk_period;
		Addr <=  "00011000110000";
		Trees_din <= x"15009c08";
		wait for Clk_period;
		Addr <=  "00011000110001";
		Trees_din <= x"15008f04";
		wait for Clk_period;
		Addr <=  "00011000110010";
		Trees_din <= x"001b18f5";
		wait for Clk_period;
		Addr <=  "00011000110011";
		Trees_din <= x"ffd918f5";
		wait for Clk_period;
		Addr <=  "00011000110100";
		Trees_din <= x"0bf98004";
		wait for Clk_period;
		Addr <=  "00011000110101";
		Trees_din <= x"ffc118f5";
		wait for Clk_period;
		Addr <=  "00011000110110";
		Trees_din <= x"004418f5";
		wait for Clk_period;
		Addr <=  "00011000110111";
		Trees_din <= x"1a00d304";
		wait for Clk_period;
		Addr <=  "00011000111000";
		Trees_din <= x"005f18f5";
		wait for Clk_period;
		Addr <=  "00011000111001";
		Trees_din <= x"ffff18f5";
		wait for Clk_period;
		Addr <=  "00011000111010";
		Trees_din <= x"14008f04";
		wait for Clk_period;
		Addr <=  "00011000111011";
		Trees_din <= x"fffc18f5";
		wait for Clk_period;
		Addr <=  "00011000111100";
		Trees_din <= x"ff9118f5";
		wait for Clk_period;
		Addr <=  "00011000111101";
		Trees_din <= x"0406be24";
		wait for Clk_period;
		Addr <=  "00011000111110";
		Trees_din <= x"12fe6204";
		wait for Clk_period;
		Addr <=  "00011000111111";
		Trees_din <= x"ff8419e1";
		wait for Clk_period;
		Addr <=  "00011001000000";
		Trees_din <= x"1a00f51c";
		wait for Clk_period;
		Addr <=  "00011001000001";
		Trees_din <= x"1a00be10";
		wait for Clk_period;
		Addr <=  "00011001000010";
		Trees_din <= x"1e008b08";
		wait for Clk_period;
		Addr <=  "00011001000011";
		Trees_din <= x"0e041104";
		wait for Clk_period;
		Addr <=  "00011001000100";
		Trees_din <= x"ff8d19e1";
		wait for Clk_period;
		Addr <=  "00011001000101";
		Trees_din <= x"002119e1";
		wait for Clk_period;
		Addr <=  "00011001000110";
		Trees_din <= x"19007204";
		wait for Clk_period;
		Addr <=  "00011001000111";
		Trees_din <= x"ffcb19e1";
		wait for Clk_period;
		Addr <=  "00011001001000";
		Trees_din <= x"004e19e1";
		wait for Clk_period;
		Addr <=  "00011001001001";
		Trees_din <= x"010a9008";
		wait for Clk_period;
		Addr <=  "00011001001010";
		Trees_din <= x"1701ad04";
		wait for Clk_period;
		Addr <=  "00011001001011";
		Trees_din <= x"004319e1";
		wait for Clk_period;
		Addr <=  "00011001001100";
		Trees_din <= x"ffdc19e1";
		wait for Clk_period;
		Addr <=  "00011001001101";
		Trees_din <= x"ff9519e1";
		wait for Clk_period;
		Addr <=  "00011001001110";
		Trees_din <= x"ff8619e1";
		wait for Clk_period;
		Addr <=  "00011001001111";
		Trees_din <= x"16011928";
		wait for Clk_period;
		Addr <=  "00011001010000";
		Trees_din <= x"14035d10";
		wait for Clk_period;
		Addr <=  "00011001010001";
		Trees_din <= x"02025f0c";
		wait for Clk_period;
		Addr <=  "00011001010010";
		Trees_din <= x"0308a908";
		wait for Clk_period;
		Addr <=  "00011001010011";
		Trees_din <= x"0f00a604";
		wait for Clk_period;
		Addr <=  "00011001010100";
		Trees_din <= x"002819e1";
		wait for Clk_period;
		Addr <=  "00011001010101";
		Trees_din <= x"009219e1";
		wait for Clk_period;
		Addr <=  "00011001010110";
		Trees_din <= x"001419e1";
		wait for Clk_period;
		Addr <=  "00011001010111";
		Trees_din <= x"ffd419e1";
		wait for Clk_period;
		Addr <=  "00011001011000";
		Trees_din <= x"17000010";
		wait for Clk_period;
		Addr <=  "00011001011001";
		Trees_din <= x"0e01e308";
		wait for Clk_period;
		Addr <=  "00011001011010";
		Trees_din <= x"0ef98b04";
		wait for Clk_period;
		Addr <=  "00011001011011";
		Trees_din <= x"ffc819e1";
		wait for Clk_period;
		Addr <=  "00011001011100";
		Trees_din <= x"005419e1";
		wait for Clk_period;
		Addr <=  "00011001011101";
		Trees_din <= x"00fcaf04";
		wait for Clk_period;
		Addr <=  "00011001011110";
		Trees_din <= x"003119e1";
		wait for Clk_period;
		Addr <=  "00011001011111";
		Trees_din <= x"ff9619e1";
		wait for Clk_period;
		Addr <=  "00011001100000";
		Trees_din <= x"13fffc04";
		wait for Clk_period;
		Addr <=  "00011001100001";
		Trees_din <= x"ff8819e1";
		wait for Clk_period;
		Addr <=  "00011001100010";
		Trees_din <= x"fff819e1";
		wait for Clk_period;
		Addr <=  "00011001100011";
		Trees_din <= x"16028714";
		wait for Clk_period;
		Addr <=  "00011001100100";
		Trees_din <= x"0b04740c";
		wait for Clk_period;
		Addr <=  "00011001100101";
		Trees_din <= x"19008d04";
		wait for Clk_period;
		Addr <=  "00011001100110";
		Trees_din <= x"000919e1";
		wait for Clk_period;
		Addr <=  "00011001100111";
		Trees_din <= x"1b003c04";
		wait for Clk_period;
		Addr <=  "00011001101000";
		Trees_din <= x"ff6e19e1";
		wait for Clk_period;
		Addr <=  "00011001101001";
		Trees_din <= x"ffe419e1";
		wait for Clk_period;
		Addr <=  "00011001101010";
		Trees_din <= x"16018d04";
		wait for Clk_period;
		Addr <=  "00011001101011";
		Trees_din <= x"ffcf19e1";
		wait for Clk_period;
		Addr <=  "00011001101100";
		Trees_din <= x"007019e1";
		wait for Clk_period;
		Addr <=  "00011001101101";
		Trees_din <= x"030a7410";
		wait for Clk_period;
		Addr <=  "00011001101110";
		Trees_din <= x"19008a08";
		wait for Clk_period;
		Addr <=  "00011001101111";
		Trees_din <= x"18004c04";
		wait for Clk_period;
		Addr <=  "00011001110000";
		Trees_din <= x"008719e1";
		wait for Clk_period;
		Addr <=  "00011001110001";
		Trees_din <= x"fffd19e1";
		wait for Clk_period;
		Addr <=  "00011001110010";
		Trees_din <= x"1a00e404";
		wait for Clk_period;
		Addr <=  "00011001110011";
		Trees_din <= x"ffe919e1";
		wait for Clk_period;
		Addr <=  "00011001110100";
		Trees_din <= x"005119e1";
		wait for Clk_period;
		Addr <=  "00011001110101";
		Trees_din <= x"14007d04";
		wait for Clk_period;
		Addr <=  "00011001110110";
		Trees_din <= x"000419e1";
		wait for Clk_period;
		Addr <=  "00011001110111";
		Trees_din <= x"ff9a19e1";
		wait for Clk_period;
		Addr <=  "00011001111000";
		Trees_din <= x"0009744c";
		wait for Clk_period;
		Addr <=  "00011001111001";
		Trees_din <= x"05fe7034";
		wait for Clk_period;
		Addr <=  "00011001111010";
		Trees_din <= x"04065f14";
		wait for Clk_period;
		Addr <=  "00011001111011";
		Trees_din <= x"17016010";
		wait for Clk_period;
		Addr <=  "00011001111100";
		Trees_din <= x"17009e08";
		wait for Clk_period;
		Addr <=  "00011001111101";
		Trees_din <= x"11045104";
		wait for Clk_period;
		Addr <=  "00011001111110";
		Trees_din <= x"ffc71a8d";
		wait for Clk_period;
		Addr <=  "00011001111111";
		Trees_din <= x"003c1a8d";
		wait for Clk_period;
		Addr <=  "00011010000000";
		Trees_din <= x"11026604";
		wait for Clk_period;
		Addr <=  "00011010000001";
		Trees_din <= x"00731a8d";
		wait for Clk_period;
		Addr <=  "00011010000010";
		Trees_din <= x"ffce1a8d";
		wait for Clk_period;
		Addr <=  "00011010000011";
		Trees_din <= x"ff7a1a8d";
		wait for Clk_period;
		Addr <=  "00011010000100";
		Trees_din <= x"0d034510";
		wait for Clk_period;
		Addr <=  "00011010000101";
		Trees_din <= x"0d02e108";
		wait for Clk_period;
		Addr <=  "00011010000110";
		Trees_din <= x"18003c04";
		wait for Clk_period;
		Addr <=  "00011010000111";
		Trees_din <= x"00371a8d";
		wait for Clk_period;
		Addr <=  "00011010001000";
		Trees_din <= x"fff81a8d";
		wait for Clk_period;
		Addr <=  "00011010001001";
		Trees_din <= x"12003304";
		wait for Clk_period;
		Addr <=  "00011010001010";
		Trees_din <= x"00231a8d";
		wait for Clk_period;
		Addr <=  "00011010001011";
		Trees_din <= x"ff801a8d";
		wait for Clk_period;
		Addr <=  "00011010001100";
		Trees_din <= x"00fb4e08";
		wait for Clk_period;
		Addr <=  "00011010001101";
		Trees_din <= x"17002d04";
		wait for Clk_period;
		Addr <=  "00011010001110";
		Trees_din <= x"001b1a8d";
		wait for Clk_period;
		Addr <=  "00011010001111";
		Trees_din <= x"ffc71a8d";
		wait for Clk_period;
		Addr <=  "00011010010000";
		Trees_din <= x"06f2f004";
		wait for Clk_period;
		Addr <=  "00011010010001";
		Trees_din <= x"ffee1a8d";
		wait for Clk_period;
		Addr <=  "00011010010010";
		Trees_din <= x"00731a8d";
		wait for Clk_period;
		Addr <=  "00011010010011";
		Trees_din <= x"0a028614";
		wait for Clk_period;
		Addr <=  "00011010010100";
		Trees_din <= x"1400c508";
		wait for Clk_period;
		Addr <=  "00011010010101";
		Trees_din <= x"15009e04";
		wait for Clk_period;
		Addr <=  "00011010010110";
		Trees_din <= x"ff951a8d";
		wait for Clk_period;
		Addr <=  "00011010010111";
		Trees_din <= x"00241a8d";
		wait for Clk_period;
		Addr <=  "00011010011000";
		Trees_din <= x"0f033208";
		wait for Clk_period;
		Addr <=  "00011010011001";
		Trees_din <= x"0c02a404";
		wait for Clk_period;
		Addr <=  "00011010011010";
		Trees_din <= x"00961a8d";
		wait for Clk_period;
		Addr <=  "00011010011011";
		Trees_din <= x"002d1a8d";
		wait for Clk_period;
		Addr <=  "00011010011100";
		Trees_din <= x"ffe11a8d";
		wait for Clk_period;
		Addr <=  "00011010011101";
		Trees_din <= x"ffb41a8d";
		wait for Clk_period;
		Addr <=  "00011010011110";
		Trees_din <= x"1d003d08";
		wait for Clk_period;
		Addr <=  "00011010011111";
		Trees_din <= x"1b003304";
		wait for Clk_period;
		Addr <=  "00011010100000";
		Trees_din <= x"ffe71a8d";
		wait for Clk_period;
		Addr <=  "00011010100001";
		Trees_din <= x"003b1a8d";
		wait for Clk_period;
		Addr <=  "00011010100010";
		Trees_din <= x"ff8a1a8d";
		wait for Clk_period;
		Addr <=  "00011010100011";
		Trees_din <= x"040a4a3c";
		wait for Clk_period;
		Addr <=  "00011010100100";
		Trees_din <= x"1d00380c";
		wait for Clk_period;
		Addr <=  "00011010100101";
		Trees_din <= x"0302da04";
		wait for Clk_period;
		Addr <=  "00011010100110";
		Trees_din <= x"ff6f1b59";
		wait for Clk_period;
		Addr <=  "00011010100111";
		Trees_din <= x"0bfaaf04";
		wait for Clk_period;
		Addr <=  "00011010101000";
		Trees_din <= x"00501b59";
		wait for Clk_period;
		Addr <=  "00011010101001";
		Trees_din <= x"ffc41b59";
		wait for Clk_period;
		Addr <=  "00011010101010";
		Trees_din <= x"1c002c14";
		wait for Clk_period;
		Addr <=  "00011010101011";
		Trees_din <= x"0801f40c";
		wait for Clk_period;
		Addr <=  "00011010101100";
		Trees_din <= x"03054208";
		wait for Clk_period;
		Addr <=  "00011010101101";
		Trees_din <= x"1703a404";
		wait for Clk_period;
		Addr <=  "00011010101110";
		Trees_din <= x"00731b59";
		wait for Clk_period;
		Addr <=  "00011010101111";
		Trees_din <= x"fffa1b59";
		wait for Clk_period;
		Addr <=  "00011010110000";
		Trees_din <= x"fff01b59";
		wait for Clk_period;
		Addr <=  "00011010110001";
		Trees_din <= x"0c024104";
		wait for Clk_period;
		Addr <=  "00011010110010";
		Trees_din <= x"00111b59";
		wait for Clk_period;
		Addr <=  "00011010110011";
		Trees_din <= x"ffa51b59";
		wait for Clk_period;
		Addr <=  "00011010110100";
		Trees_din <= x"1c002e0c";
		wait for Clk_period;
		Addr <=  "00011010110101";
		Trees_din <= x"0efcb004";
		wait for Clk_period;
		Addr <=  "00011010110110";
		Trees_din <= x"00281b59";
		wait for Clk_period;
		Addr <=  "00011010110111";
		Trees_din <= x"14022404";
		wait for Clk_period;
		Addr <=  "00011010111000";
		Trees_din <= x"ff701b59";
		wait for Clk_period;
		Addr <=  "00011010111001";
		Trees_din <= x"ffe61b59";
		wait for Clk_period;
		Addr <=  "00011010111010";
		Trees_din <= x"1c003508";
		wait for Clk_period;
		Addr <=  "00011010111011";
		Trees_din <= x"05fd4604";
		wait for Clk_period;
		Addr <=  "00011010111100";
		Trees_din <= x"ffea1b59";
		wait for Clk_period;
		Addr <=  "00011010111101";
		Trees_din <= x"005b1b59";
		wait for Clk_period;
		Addr <=  "00011010111110";
		Trees_din <= x"00046404";
		wait for Clk_period;
		Addr <=  "00011010111111";
		Trees_din <= x"fff71b59";
		wait for Clk_period;
		Addr <=  "00011011000000";
		Trees_din <= x"ffa71b59";
		wait for Clk_period;
		Addr <=  "00011011000001";
		Trees_din <= x"00feb724";
		wait for Clk_period;
		Addr <=  "00011011000010";
		Trees_din <= x"0b028214";
		wait for Clk_period;
		Addr <=  "00011011000011";
		Trees_din <= x"1e00700c";
		wait for Clk_period;
		Addr <=  "00011011000100";
		Trees_din <= x"14012704";
		wait for Clk_period;
		Addr <=  "00011011000101";
		Trees_din <= x"00071b59";
		wait for Clk_period;
		Addr <=  "00011011000110";
		Trees_din <= x"02ff2a04";
		wait for Clk_period;
		Addr <=  "00011011000111";
		Trees_din <= x"fff61b59";
		wait for Clk_period;
		Addr <=  "00011011001000";
		Trees_din <= x"ff851b59";
		wait for Clk_period;
		Addr <=  "00011011001001";
		Trees_din <= x"07005804";
		wait for Clk_period;
		Addr <=  "00011011001010";
		Trees_din <= x"005b1b59";
		wait for Clk_period;
		Addr <=  "00011011001011";
		Trees_din <= x"ffe61b59";
		wait for Clk_period;
		Addr <=  "00011011001100";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00011011001101";
		Trees_din <= x"00691b59";
		wait for Clk_period;
		Addr <=  "00011011001110";
		Trees_din <= x"18004a08";
		wait for Clk_period;
		Addr <=  "00011011001111";
		Trees_din <= x"0101fc04";
		wait for Clk_period;
		Addr <=  "00011011010000";
		Trees_din <= x"ffa71b59";
		wait for Clk_period;
		Addr <=  "00011011010001";
		Trees_din <= x"fffc1b59";
		wait for Clk_period;
		Addr <=  "00011011010010";
		Trees_din <= x"00451b59";
		wait for Clk_period;
		Addr <=  "00011011010011";
		Trees_din <= x"0106e504";
		wait for Clk_period;
		Addr <=  "00011011010100";
		Trees_din <= x"00841b59";
		wait for Clk_period;
		Addr <=  "00011011010101";
		Trees_din <= x"ffee1b59";
		wait for Clk_period;
		Addr <=  "00011011010110";
		Trees_din <= x"04faa904";
		wait for Clk_period;
		Addr <=  "00011011010111";
		Trees_din <= x"ffa11c1d";
		wait for Clk_period;
		Addr <=  "00011011011000";
		Trees_din <= x"1900a83c";
		wait for Clk_period;
		Addr <=  "00011011011001";
		Trees_din <= x"0700581c";
		wait for Clk_period;
		Addr <=  "00011011011010";
		Trees_din <= x"1603c910";
		wait for Clk_period;
		Addr <=  "00011011011011";
		Trees_din <= x"1c003608";
		wait for Clk_period;
		Addr <=  "00011011011100";
		Trees_din <= x"09005404";
		wait for Clk_period;
		Addr <=  "00011011011101";
		Trees_din <= x"000a1c1d";
		wait for Clk_period;
		Addr <=  "00011011011110";
		Trees_din <= x"00701c1d";
		wait for Clk_period;
		Addr <=  "00011011011111";
		Trees_din <= x"0a028704";
		wait for Clk_period;
		Addr <=  "00011011100000";
		Trees_din <= x"001a1c1d";
		wait for Clk_period;
		Addr <=  "00011011100001";
		Trees_din <= x"ffbd1c1d";
		wait for Clk_period;
		Addr <=  "00011011100010";
		Trees_din <= x"04077804";
		wait for Clk_period;
		Addr <=  "00011011100011";
		Trees_din <= x"ff901c1d";
		wait for Clk_period;
		Addr <=  "00011011100100";
		Trees_din <= x"11011304";
		wait for Clk_period;
		Addr <=  "00011011100101";
		Trees_din <= x"ffd21c1d";
		wait for Clk_period;
		Addr <=  "00011011100110";
		Trees_din <= x"00541c1d";
		wait for Clk_period;
		Addr <=  "00011011100111";
		Trees_din <= x"11012610";
		wait for Clk_period;
		Addr <=  "00011011101000";
		Trees_din <= x"20040008";
		wait for Clk_period;
		Addr <=  "00011011101001";
		Trees_din <= x"1b003b04";
		wait for Clk_period;
		Addr <=  "00011011101010";
		Trees_din <= x"fff41c1d";
		wait for Clk_period;
		Addr <=  "00011011101011";
		Trees_din <= x"00821c1d";
		wait for Clk_period;
		Addr <=  "00011011101100";
		Trees_din <= x"19009004";
		wait for Clk_period;
		Addr <=  "00011011101101";
		Trees_din <= x"003a1c1d";
		wait for Clk_period;
		Addr <=  "00011011101110";
		Trees_din <= x"ffad1c1d";
		wait for Clk_period;
		Addr <=  "00011011101111";
		Trees_din <= x"06f7d508";
		wait for Clk_period;
		Addr <=  "00011011110000";
		Trees_din <= x"1104d504";
		wait for Clk_period;
		Addr <=  "00011011110001";
		Trees_din <= x"ffab1c1d";
		wait for Clk_period;
		Addr <=  "00011011110010";
		Trees_din <= x"00491c1d";
		wait for Clk_period;
		Addr <=  "00011011110011";
		Trees_din <= x"1a00bc04";
		wait for Clk_period;
		Addr <=  "00011011110100";
		Trees_din <= x"ffa81c1d";
		wait for Clk_period;
		Addr <=  "00011011110101";
		Trees_din <= x"00771c1d";
		wait for Clk_period;
		Addr <=  "00011011110110";
		Trees_din <= x"1c002a18";
		wait for Clk_period;
		Addr <=  "00011011110111";
		Trees_din <= x"1c002508";
		wait for Clk_period;
		Addr <=  "00011011111000";
		Trees_din <= x"01034104";
		wait for Clk_period;
		Addr <=  "00011011111001";
		Trees_din <= x"fffe1c1d";
		wait for Clk_period;
		Addr <=  "00011011111010";
		Trees_din <= x"ff9d1c1d";
		wait for Clk_period;
		Addr <=  "00011011111011";
		Trees_din <= x"04060d08";
		wait for Clk_period;
		Addr <=  "00011011111100";
		Trees_din <= x"05fdfd04";
		wait for Clk_period;
		Addr <=  "00011011111101";
		Trees_din <= x"ffb11c1d";
		wait for Clk_period;
		Addr <=  "00011011111110";
		Trees_din <= x"00041c1d";
		wait for Clk_period;
		Addr <=  "00011011111111";
		Trees_din <= x"00001404";
		wait for Clk_period;
		Addr <=  "00011100000000";
		Trees_din <= x"007a1c1d";
		wait for Clk_period;
		Addr <=  "00011100000001";
		Trees_din <= x"00141c1d";
		wait for Clk_period;
		Addr <=  "00011100000010";
		Trees_din <= x"01031d08";
		wait for Clk_period;
		Addr <=  "00011100000011";
		Trees_din <= x"0d015f04";
		wait for Clk_period;
		Addr <=  "00011100000100";
		Trees_din <= x"00321c1d";
		wait for Clk_period;
		Addr <=  "00011100000101";
		Trees_din <= x"ffba1c1d";
		wait for Clk_period;
		Addr <=  "00011100000110";
		Trees_din <= x"ff721c1d";
		wait for Clk_period;
		Addr <=  "00011100000111";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00011100001000";
		Trees_din <= x"040a4a3c";
		wait for Clk_period;
		Addr <=  "00011100001001";
		Trees_din <= x"1d00380c";
		wait for Clk_period;
		Addr <=  "00011100001010";
		Trees_din <= x"0302da04";
		wait for Clk_period;
		Addr <=  "00011100001011";
		Trees_din <= x"ff791cf5";
		wait for Clk_period;
		Addr <=  "00011100001100";
		Trees_din <= x"0bfaaf04";
		wait for Clk_period;
		Addr <=  "00011100001101";
		Trees_din <= x"004b1cf5";
		wait for Clk_period;
		Addr <=  "00011100001110";
		Trees_din <= x"ffc71cf5";
		wait for Clk_period;
		Addr <=  "00011100001111";
		Trees_din <= x"1c002c14";
		wait for Clk_period;
		Addr <=  "00011100010000";
		Trees_din <= x"0801f40c";
		wait for Clk_period;
		Addr <=  "00011100010001";
		Trees_din <= x"03054208";
		wait for Clk_period;
		Addr <=  "00011100010010";
		Trees_din <= x"0401dd04";
		wait for Clk_period;
		Addr <=  "00011100010011";
		Trees_din <= x"00021cf5";
		wait for Clk_period;
		Addr <=  "00011100010100";
		Trees_din <= x"00691cf5";
		wait for Clk_period;
		Addr <=  "00011100010101";
		Trees_din <= x"fff11cf5";
		wait for Clk_period;
		Addr <=  "00011100010110";
		Trees_din <= x"0c024104";
		wait for Clk_period;
		Addr <=  "00011100010111";
		Trees_din <= x"000f1cf5";
		wait for Clk_period;
		Addr <=  "00011100011000";
		Trees_din <= x"ffad1cf5";
		wait for Clk_period;
		Addr <=  "00011100011001";
		Trees_din <= x"1c002e0c";
		wait for Clk_period;
		Addr <=  "00011100011010";
		Trees_din <= x"0efcb004";
		wait for Clk_period;
		Addr <=  "00011100011011";
		Trees_din <= x"00231cf5";
		wait for Clk_period;
		Addr <=  "00011100011100";
		Trees_din <= x"14022404";
		wait for Clk_period;
		Addr <=  "00011100011101";
		Trees_din <= x"ff781cf5";
		wait for Clk_period;
		Addr <=  "00011100011110";
		Trees_din <= x"ffe71cf5";
		wait for Clk_period;
		Addr <=  "00011100011111";
		Trees_din <= x"05fa9208";
		wait for Clk_period;
		Addr <=  "00011100100000";
		Trees_din <= x"0d03bf04";
		wait for Clk_period;
		Addr <=  "00011100100001";
		Trees_din <= x"ffaf1cf5";
		wait for Clk_period;
		Addr <=  "00011100100010";
		Trees_din <= x"00291cf5";
		wait for Clk_period;
		Addr <=  "00011100100011";
		Trees_din <= x"15009e04";
		wait for Clk_period;
		Addr <=  "00011100100100";
		Trees_din <= x"fff81cf5";
		wait for Clk_period;
		Addr <=  "00011100100101";
		Trees_din <= x"004c1cf5";
		wait for Clk_period;
		Addr <=  "00011100100110";
		Trees_din <= x"030a7428";
		wait for Clk_period;
		Addr <=  "00011100100111";
		Trees_din <= x"01068718";
		wait for Clk_period;
		Addr <=  "00011100101000";
		Trees_din <= x"0900570c";
		wait for Clk_period;
		Addr <=  "00011100101001";
		Trees_din <= x"07005b08";
		wait for Clk_period;
		Addr <=  "00011100101010";
		Trees_din <= x"1202c604";
		wait for Clk_period;
		Addr <=  "00011100101011";
		Trees_din <= x"007d1cf5";
		wait for Clk_period;
		Addr <=  "00011100101100";
		Trees_din <= x"001f1cf5";
		wait for Clk_period;
		Addr <=  "00011100101101";
		Trees_din <= x"00101cf5";
		wait for Clk_period;
		Addr <=  "00011100101110";
		Trees_din <= x"06f34c04";
		wait for Clk_period;
		Addr <=  "00011100101111";
		Trees_din <= x"003e1cf5";
		wait for Clk_period;
		Addr <=  "00011100110000";
		Trees_din <= x"1c003a04";
		wait for Clk_period;
		Addr <=  "00011100110001";
		Trees_din <= x"00051cf5";
		wait for Clk_period;
		Addr <=  "00011100110010";
		Trees_din <= x"ffb11cf5";
		wait for Clk_period;
		Addr <=  "00011100110011";
		Trees_din <= x"13ffe60c";
		wait for Clk_period;
		Addr <=  "00011100110100";
		Trees_din <= x"040c1204";
		wait for Clk_period;
		Addr <=  "00011100110101";
		Trees_din <= x"ff981cf5";
		wait for Clk_period;
		Addr <=  "00011100110110";
		Trees_din <= x"1a00d204";
		wait for Clk_period;
		Addr <=  "00011100110111";
		Trees_din <= x"004c1cf5";
		wait for Clk_period;
		Addr <=  "00011100111000";
		Trees_din <= x"ffcd1cf5";
		wait for Clk_period;
		Addr <=  "00011100111001";
		Trees_din <= x"005e1cf5";
		wait for Clk_period;
		Addr <=  "00011100111010";
		Trees_din <= x"0f00a604";
		wait for Clk_period;
		Addr <=  "00011100111011";
		Trees_din <= x"00071cf5";
		wait for Clk_period;
		Addr <=  "00011100111100";
		Trees_din <= x"ffa91cf5";
		wait for Clk_period;
		Addr <=  "00011100111101";
		Trees_din <= x"00097434";
		wait for Clk_period;
		Addr <=  "00011100111110";
		Trees_din <= x"1e008b24";
		wait for Clk_period;
		Addr <=  "00011100111111";
		Trees_din <= x"18004c18";
		wait for Clk_period;
		Addr <=  "00011101000000";
		Trees_din <= x"09005b10";
		wait for Clk_period;
		Addr <=  "00011101000001";
		Trees_din <= x"0c006108";
		wait for Clk_period;
		Addr <=  "00011101000010";
		Trees_din <= x"0b042604";
		wait for Clk_period;
		Addr <=  "00011101000011";
		Trees_din <= x"004e1d69";
		wait for Clk_period;
		Addr <=  "00011101000100";
		Trees_din <= x"ffe11d69";
		wait for Clk_period;
		Addr <=  "00011101000101";
		Trees_din <= x"0c021f04";
		wait for Clk_period;
		Addr <=  "00011101000110";
		Trees_din <= x"ffde1d69";
		wait for Clk_period;
		Addr <=  "00011101000111";
		Trees_din <= x"00101d69";
		wait for Clk_period;
		Addr <=  "00011101001000";
		Trees_din <= x"1900a004";
		wait for Clk_period;
		Addr <=  "00011101001001";
		Trees_din <= x"00001d69";
		wait for Clk_period;
		Addr <=  "00011101001010";
		Trees_din <= x"00791d69";
		wait for Clk_period;
		Addr <=  "00011101001011";
		Trees_din <= x"0408ca04";
		wait for Clk_period;
		Addr <=  "00011101001100";
		Trees_din <= x"ff901d69";
		wait for Clk_period;
		Addr <=  "00011101001101";
		Trees_din <= x"1200e704";
		wait for Clk_period;
		Addr <=  "00011101001110";
		Trees_din <= x"00221d69";
		wait for Clk_period;
		Addr <=  "00011101001111";
		Trees_din <= x"ffe91d69";
		wait for Clk_period;
		Addr <=  "00011101010000";
		Trees_din <= x"19007204";
		wait for Clk_period;
		Addr <=  "00011101010001";
		Trees_din <= x"ffc41d69";
		wait for Clk_period;
		Addr <=  "00011101010010";
		Trees_din <= x"15007b08";
		wait for Clk_period;
		Addr <=  "00011101010011";
		Trees_din <= x"08005004";
		wait for Clk_period;
		Addr <=  "00011101010100";
		Trees_din <= x"ffee1d69";
		wait for Clk_period;
		Addr <=  "00011101010101";
		Trees_din <= x"00261d69";
		wait for Clk_period;
		Addr <=  "00011101010110";
		Trees_din <= x"007f1d69";
		wait for Clk_period;
		Addr <=  "00011101010111";
		Trees_din <= x"1d003d04";
		wait for Clk_period;
		Addr <=  "00011101011000";
		Trees_din <= x"000f1d69";
		wait for Clk_period;
		Addr <=  "00011101011001";
		Trees_din <= x"ff931d69";
		wait for Clk_period;
		Addr <=  "00011101011010";
		Trees_din <= x"040a4a38";
		wait for Clk_period;
		Addr <=  "00011101011011";
		Trees_din <= x"1d00380c";
		wait for Clk_period;
		Addr <=  "00011101011100";
		Trees_din <= x"0302da04";
		wait for Clk_period;
		Addr <=  "00011101011101";
		Trees_din <= x"ff7f1e2d";
		wait for Clk_period;
		Addr <=  "00011101011110";
		Trees_din <= x"0bfaaf04";
		wait for Clk_period;
		Addr <=  "00011101011111";
		Trees_din <= x"00451e2d";
		wait for Clk_period;
		Addr <=  "00011101100000";
		Trees_din <= x"ffcd1e2d";
		wait for Clk_period;
		Addr <=  "00011101100001";
		Trees_din <= x"1c002c18";
		wait for Clk_period;
		Addr <=  "00011101100010";
		Trees_din <= x"02012d10";
		wait for Clk_period;
		Addr <=  "00011101100011";
		Trees_din <= x"10040608";
		wait for Clk_period;
		Addr <=  "00011101100100";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00011101100101";
		Trees_din <= x"00051e2d";
		wait for Clk_period;
		Addr <=  "00011101100110";
		Trees_din <= x"00771e2d";
		wait for Clk_period;
		Addr <=  "00011101100111";
		Trees_din <= x"06f73504";
		wait for Clk_period;
		Addr <=  "00011101101000";
		Trees_din <= x"ffc81e2d";
		wait for Clk_period;
		Addr <=  "00011101101001";
		Trees_din <= x"00421e2d";
		wait for Clk_period;
		Addr <=  "00011101101010";
		Trees_din <= x"02045404";
		wait for Clk_period;
		Addr <=  "00011101101011";
		Trees_din <= x"ffbd1e2d";
		wait for Clk_period;
		Addr <=  "00011101101100";
		Trees_din <= x"00071e2d";
		wait for Clk_period;
		Addr <=  "00011101101101";
		Trees_din <= x"010c6810";
		wait for Clk_period;
		Addr <=  "00011101101110";
		Trees_din <= x"00fa9208";
		wait for Clk_period;
		Addr <=  "00011101101111";
		Trees_din <= x"0c029704";
		wait for Clk_period;
		Addr <=  "00011101110000";
		Trees_din <= x"ff941e2d";
		wait for Clk_period;
		Addr <=  "00011101110001";
		Trees_din <= x"00131e2d";
		wait for Clk_period;
		Addr <=  "00011101110010";
		Trees_din <= x"00fd2504";
		wait for Clk_period;
		Addr <=  "00011101110011";
		Trees_din <= x"00431e2d";
		wait for Clk_period;
		Addr <=  "00011101110100";
		Trees_din <= x"fff11e2d";
		wait for Clk_period;
		Addr <=  "00011101110101";
		Trees_din <= x"ff991e2d";
		wait for Clk_period;
		Addr <=  "00011101110110";
		Trees_din <= x"00feb724";
		wait for Clk_period;
		Addr <=  "00011101110111";
		Trees_din <= x"0b028214";
		wait for Clk_period;
		Addr <=  "00011101111000";
		Trees_din <= x"1e00700c";
		wait for Clk_period;
		Addr <=  "00011101111001";
		Trees_din <= x"14012704";
		wait for Clk_period;
		Addr <=  "00011101111010";
		Trees_din <= x"00071e2d";
		wait for Clk_period;
		Addr <=  "00011101111011";
		Trees_din <= x"02ff2a04";
		wait for Clk_period;
		Addr <=  "00011101111100";
		Trees_din <= x"fffd1e2d";
		wait for Clk_period;
		Addr <=  "00011101111101";
		Trees_din <= x"ff911e2d";
		wait for Clk_period;
		Addr <=  "00011101111110";
		Trees_din <= x"13ffeb04";
		wait for Clk_period;
		Addr <=  "00011101111111";
		Trees_din <= x"fff61e2d";
		wait for Clk_period;
		Addr <=  "00011110000000";
		Trees_din <= x"00451e2d";
		wait for Clk_period;
		Addr <=  "00011110000001";
		Trees_din <= x"07005908";
		wait for Clk_period;
		Addr <=  "00011110000010";
		Trees_din <= x"0f00f204";
		wait for Clk_period;
		Addr <=  "00011110000011";
		Trees_din <= x"006c1e2d";
		wait for Clk_period;
		Addr <=  "00011110000100";
		Trees_din <= x"001e1e2d";
		wait for Clk_period;
		Addr <=  "00011110000101";
		Trees_din <= x"17000004";
		wait for Clk_period;
		Addr <=  "00011110000110";
		Trees_din <= x"002d1e2d";
		wait for Clk_period;
		Addr <=  "00011110000111";
		Trees_din <= x"ffc21e2d";
		wait for Clk_period;
		Addr <=  "00011110001000";
		Trees_din <= x"0106e504";
		wait for Clk_period;
		Addr <=  "00011110001001";
		Trees_din <= x"00791e2d";
		wait for Clk_period;
		Addr <=  "00011110001010";
		Trees_din <= x"fff11e2d";
		wait for Clk_period;
		Addr <=  "00011110001011";
		Trees_din <= x"040e643c";
		wait for Clk_period;
		Addr <=  "00011110001100";
		Trees_din <= x"03fb1e08";
		wait for Clk_period;
		Addr <=  "00011110001101";
		Trees_din <= x"01031d04";
		wait for Clk_period;
		Addr <=  "00011110001110";
		Trees_din <= x"00171eb1";
		wait for Clk_period;
		Addr <=  "00011110001111";
		Trees_din <= x"ff961eb1";
		wait for Clk_period;
		Addr <=  "00011110010000";
		Trees_din <= x"1603c91c";
		wait for Clk_period;
		Addr <=  "00011110010001";
		Trees_din <= x"1900a810";
		wait for Clk_period;
		Addr <=  "00011110010010";
		Trees_din <= x"07005608";
		wait for Clk_period;
		Addr <=  "00011110010011";
		Trees_din <= x"19009b04";
		wait for Clk_period;
		Addr <=  "00011110010100";
		Trees_din <= x"00031eb1";
		wait for Clk_period;
		Addr <=  "00011110010101";
		Trees_din <= x"00541eb1";
		wait for Clk_period;
		Addr <=  "00011110010110";
		Trees_din <= x"0c006e04";
		wait for Clk_period;
		Addr <=  "00011110010111";
		Trees_din <= x"00461eb1";
		wait for Clk_period;
		Addr <=  "00011110011000";
		Trees_din <= x"ffea1eb1";
		wait for Clk_period;
		Addr <=  "00011110011001";
		Trees_din <= x"1900aa04";
		wait for Clk_period;
		Addr <=  "00011110011010";
		Trees_din <= x"ff931eb1";
		wait for Clk_period;
		Addr <=  "00011110011011";
		Trees_din <= x"02ff7304";
		wait for Clk_period;
		Addr <=  "00011110011100";
		Trees_din <= x"00321eb1";
		wait for Clk_period;
		Addr <=  "00011110011101";
		Trees_din <= x"ffc41eb1";
		wait for Clk_period;
		Addr <=  "00011110011110";
		Trees_din <= x"04070608";
		wait for Clk_period;
		Addr <=  "00011110011111";
		Trees_din <= x"1900a604";
		wait for Clk_period;
		Addr <=  "00011110100000";
		Trees_din <= x"ff7e1eb1";
		wait for Clk_period;
		Addr <=  "00011110100001";
		Trees_din <= x"001e1eb1";
		wait for Clk_period;
		Addr <=  "00011110100010";
		Trees_din <= x"1200a408";
		wait for Clk_period;
		Addr <=  "00011110100011";
		Trees_din <= x"00fcaf04";
		wait for Clk_period;
		Addr <=  "00011110100100";
		Trees_din <= x"001e1eb1";
		wait for Clk_period;
		Addr <=  "00011110100101";
		Trees_din <= x"ffa21eb1";
		wait for Clk_period;
		Addr <=  "00011110100110";
		Trees_din <= x"17034504";
		wait for Clk_period;
		Addr <=  "00011110100111";
		Trees_din <= x"fff21eb1";
		wait for Clk_period;
		Addr <=  "00011110101000";
		Trees_din <= x"00621eb1";
		wait for Clk_period;
		Addr <=  "00011110101001";
		Trees_din <= x"1a00d304";
		wait for Clk_period;
		Addr <=  "00011110101010";
		Trees_din <= x"00551eb1";
		wait for Clk_period;
		Addr <=  "00011110101011";
		Trees_din <= x"00001eb1";
		wait for Clk_period;
		Addr <=  "00011110101100";
		Trees_din <= x"040c1228";
		wait for Clk_period;
		Addr <=  "00011110101101";
		Trees_din <= x"07004a04";
		wait for Clk_period;
		Addr <=  "00011110101110";
		Trees_din <= x"ffac1f1d";
		wait for Clk_period;
		Addr <=  "00011110101111";
		Trees_din <= x"03fb1e08";
		wait for Clk_period;
		Addr <=  "00011110110000";
		Trees_din <= x"0afb1304";
		wait for Clk_period;
		Addr <=  "00011110110001";
		Trees_din <= x"fffb1f1d";
		wait for Clk_period;
		Addr <=  "00011110110010";
		Trees_din <= x"ff9e1f1d";
		wait for Clk_period;
		Addr <=  "00011110110011";
		Trees_din <= x"0e045b10";
		wait for Clk_period;
		Addr <=  "00011110110100";
		Trees_din <= x"06f3d608";
		wait for Clk_period;
		Addr <=  "00011110110101";
		Trees_din <= x"0afccf04";
		wait for Clk_period;
		Addr <=  "00011110110110";
		Trees_din <= x"000a1f1d";
		wait for Clk_period;
		Addr <=  "00011110110111";
		Trees_din <= x"ffad1f1d";
		wait for Clk_period;
		Addr <=  "00011110111000";
		Trees_din <= x"1d003804";
		wait for Clk_period;
		Addr <=  "00011110111001";
		Trees_din <= x"ffb21f1d";
		wait for Clk_period;
		Addr <=  "00011110111010";
		Trees_din <= x"000c1f1d";
		wait for Clk_period;
		Addr <=  "00011110111011";
		Trees_din <= x"1401d304";
		wait for Clk_period;
		Addr <=  "00011110111100";
		Trees_din <= x"ffda1f1d";
		wait for Clk_period;
		Addr <=  "00011110111101";
		Trees_din <= x"0f02ce04";
		wait for Clk_period;
		Addr <=  "00011110111110";
		Trees_din <= x"00751f1d";
		wait for Clk_period;
		Addr <=  "00011110111111";
		Trees_din <= x"00071f1d";
		wait for Clk_period;
		Addr <=  "00011111000000";
		Trees_din <= x"030a740c";
		wait for Clk_period;
		Addr <=  "00011111000001";
		Trees_din <= x"0202d908";
		wait for Clk_period;
		Addr <=  "00011111000010";
		Trees_din <= x"12fe6c04";
		wait for Clk_period;
		Addr <=  "00011111000011";
		Trees_din <= x"ffec1f1d";
		wait for Clk_period;
		Addr <=  "00011111000100";
		Trees_din <= x"00731f1d";
		wait for Clk_period;
		Addr <=  "00011111000101";
		Trees_din <= x"ffe61f1d";
		wait for Clk_period;
		Addr <=  "00011111000110";
		Trees_din <= x"ffd11f1d";
		wait for Clk_period;
		Addr <=  "00011111000111";
		Trees_din <= x"0406be30";
		wait for Clk_period;
		Addr <=  "00011111001000";
		Trees_din <= x"12fe6204";
		wait for Clk_period;
		Addr <=  "00011111001001";
		Trees_din <= x"ff922009";
		wait for Clk_period;
		Addr <=  "00011111001010";
		Trees_din <= x"1e005d0c";
		wait for Clk_period;
		Addr <=  "00011111001011";
		Trees_din <= x"1603e308";
		wait for Clk_period;
		Addr <=  "00011111001100";
		Trees_din <= x"05fe0504";
		wait for Clk_period;
		Addr <=  "00011111001101";
		Trees_din <= x"ff952009";
		wait for Clk_period;
		Addr <=  "00011111001110";
		Trees_din <= x"fff72009";
		wait for Clk_period;
		Addr <=  "00011111001111";
		Trees_din <= x"00152009";
		wait for Clk_period;
		Addr <=  "00011111010000";
		Trees_din <= x"1e006a10";
		wait for Clk_period;
		Addr <=  "00011111010001";
		Trees_din <= x"12011308";
		wait for Clk_period;
		Addr <=  "00011111010010";
		Trees_din <= x"1603c904";
		wait for Clk_period;
		Addr <=  "00011111010011";
		Trees_din <= x"00722009";
		wait for Clk_period;
		Addr <=  "00011111010100";
		Trees_din <= x"fffa2009";
		wait for Clk_period;
		Addr <=  "00011111010101";
		Trees_din <= x"05fdec04";
		wait for Clk_period;
		Addr <=  "00011111010110";
		Trees_din <= x"ffb52009";
		wait for Clk_period;
		Addr <=  "00011111010111";
		Trees_din <= x"00292009";
		wait for Clk_period;
		Addr <=  "00011111011000";
		Trees_din <= x"12019d08";
		wait for Clk_period;
		Addr <=  "00011111011001";
		Trees_din <= x"09005304";
		wait for Clk_period;
		Addr <=  "00011111011010";
		Trees_din <= x"ffee2009";
		wait for Clk_period;
		Addr <=  "00011111011011";
		Trees_din <= x"ff8b2009";
		wait for Clk_period;
		Addr <=  "00011111011100";
		Trees_din <= x"02007704";
		wait for Clk_period;
		Addr <=  "00011111011101";
		Trees_din <= x"ffa32009";
		wait for Clk_period;
		Addr <=  "00011111011110";
		Trees_din <= x"002f2009";
		wait for Clk_period;
		Addr <=  "00011111011111";
		Trees_din <= x"16011920";
		wait for Clk_period;
		Addr <=  "00011111100000";
		Trees_din <= x"14035d08";
		wait for Clk_period;
		Addr <=  "00011111100001";
		Trees_din <= x"0200a004";
		wait for Clk_period;
		Addr <=  "00011111100010";
		Trees_din <= x"00642009";
		wait for Clk_period;
		Addr <=  "00011111100011";
		Trees_din <= x"000c2009";
		wait for Clk_period;
		Addr <=  "00011111100100";
		Trees_din <= x"00feee10";
		wait for Clk_period;
		Addr <=  "00011111100101";
		Trees_din <= x"10028408";
		wait for Clk_period;
		Addr <=  "00011111100110";
		Trees_din <= x"05faf304";
		wait for Clk_period;
		Addr <=  "00011111100111";
		Trees_din <= x"ffcc2009";
		wait for Clk_period;
		Addr <=  "00011111101000";
		Trees_din <= x"001a2009";
		wait for Clk_period;
		Addr <=  "00011111101001";
		Trees_din <= x"0103ae04";
		wait for Clk_period;
		Addr <=  "00011111101010";
		Trees_din <= x"001e2009";
		wait for Clk_period;
		Addr <=  "00011111101011";
		Trees_din <= x"006a2009";
		wait for Clk_period;
		Addr <=  "00011111101100";
		Trees_din <= x"01036504";
		wait for Clk_period;
		Addr <=  "00011111101101";
		Trees_din <= x"00182009";
		wait for Clk_period;
		Addr <=  "00011111101110";
		Trees_din <= x"ff992009";
		wait for Clk_period;
		Addr <=  "00011111101111";
		Trees_din <= x"16028710";
		wait for Clk_period;
		Addr <=  "00011111110000";
		Trees_din <= x"0b047408";
		wait for Clk_period;
		Addr <=  "00011111110001";
		Trees_din <= x"19008d04";
		wait for Clk_period;
		Addr <=  "00011111110010";
		Trees_din <= x"00052009";
		wait for Clk_period;
		Addr <=  "00011111110011";
		Trees_din <= x"ff8d2009";
		wait for Clk_period;
		Addr <=  "00011111110100";
		Trees_din <= x"0a01c104";
		wait for Clk_period;
		Addr <=  "00011111110101";
		Trees_din <= x"ffef2009";
		wait for Clk_period;
		Addr <=  "00011111110110";
		Trees_din <= x"00592009";
		wait for Clk_period;
		Addr <=  "00011111110111";
		Trees_din <= x"030a7410";
		wait for Clk_period;
		Addr <=  "00011111111000";
		Trees_din <= x"12018b08";
		wait for Clk_period;
		Addr <=  "00011111111001";
		Trees_din <= x"0e014504";
		wait for Clk_period;
		Addr <=  "00011111111010";
		Trees_din <= x"00202009";
		wait for Clk_period;
		Addr <=  "00011111111011";
		Trees_din <= x"ffa72009";
		wait for Clk_period;
		Addr <=  "00011111111100";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00011111111101";
		Trees_din <= x"005d2009";
		wait for Clk_period;
		Addr <=  "00011111111110";
		Trees_din <= x"ffd12009";
		wait for Clk_period;
		Addr <=  "00011111111111";
		Trees_din <= x"1200fb04";
		wait for Clk_period;
		Addr <=  "00100000000000";
		Trees_din <= x"fffb2009";
		wait for Clk_period;
		Addr <=  "00100000000001";
		Trees_din <= x"ffac2009";
		wait for Clk_period;
		Addr <=  "00100000000010";
		Trees_din <= x"0404aa28";
		wait for Clk_period;
		Addr <=  "00100000000011";
		Trees_din <= x"15008d10";
		wait for Clk_period;
		Addr <=  "00100000000100";
		Trees_din <= x"12010f04";
		wait for Clk_period;
		Addr <=  "00100000000101";
		Trees_din <= x"ffab20d5";
		wait for Clk_period;
		Addr <=  "00100000000110";
		Trees_din <= x"1a00b908";
		wait for Clk_period;
		Addr <=  "00100000000111";
		Trees_din <= x"1c004b04";
		wait for Clk_period;
		Addr <=  "00100000001000";
		Trees_din <= x"ffc220d5";
		wait for Clk_period;
		Addr <=  "00100000001001";
		Trees_din <= x"004720d5";
		wait for Clk_period;
		Addr <=  "00100000001010";
		Trees_din <= x"007020d5";
		wait for Clk_period;
		Addr <=  "00100000001011";
		Trees_din <= x"15009d04";
		wait for Clk_period;
		Addr <=  "00100000001100";
		Trees_din <= x"ff8a20d5";
		wait for Clk_period;
		Addr <=  "00100000001101";
		Trees_din <= x"1500a008";
		wait for Clk_period;
		Addr <=  "00100000001110";
		Trees_din <= x"0f003b04";
		wait for Clk_period;
		Addr <=  "00100000001111";
		Trees_din <= x"005d20d5";
		wait for Clk_period;
		Addr <=  "00100000010000";
		Trees_din <= x"001320d5";
		wait for Clk_period;
		Addr <=  "00100000010001";
		Trees_din <= x"0afc5308";
		wait for Clk_period;
		Addr <=  "00100000010010";
		Trees_din <= x"06f84404";
		wait for Clk_period;
		Addr <=  "00100000010011";
		Trees_din <= x"ffe020d5";
		wait for Clk_period;
		Addr <=  "00100000010100";
		Trees_din <= x"002220d5";
		wait for Clk_period;
		Addr <=  "00100000010101";
		Trees_din <= x"ff9820d5";
		wait for Clk_period;
		Addr <=  "00100000010110";
		Trees_din <= x"0d034d2c";
		wait for Clk_period;
		Addr <=  "00100000010111";
		Trees_din <= x"0d02e120";
		wait for Clk_period;
		Addr <=  "00100000011000";
		Trees_din <= x"08014810";
		wait for Clk_period;
		Addr <=  "00100000011001";
		Trees_din <= x"04086a08";
		wait for Clk_period;
		Addr <=  "00100000011010";
		Trees_din <= x"0305c704";
		wait for Clk_period;
		Addr <=  "00100000011011";
		Trees_din <= x"ff9e20d5";
		wait for Clk_period;
		Addr <=  "00100000011100";
		Trees_din <= x"000920d5";
		wait for Clk_period;
		Addr <=  "00100000011101";
		Trees_din <= x"10f9d204";
		wait for Clk_period;
		Addr <=  "00100000011110";
		Trees_din <= x"ffb020d5";
		wait for Clk_period;
		Addr <=  "00100000011111";
		Trees_din <= x"002120d5";
		wait for Clk_period;
		Addr <=  "00100000100000";
		Trees_din <= x"0308a908";
		wait for Clk_period;
		Addr <=  "00100000100001";
		Trees_din <= x"07005b04";
		wait for Clk_period;
		Addr <=  "00100000100010";
		Trees_din <= x"003f20d5";
		wait for Clk_period;
		Addr <=  "00100000100011";
		Trees_din <= x"ffb120d5";
		wait for Clk_period;
		Addr <=  "00100000100100";
		Trees_din <= x"0c023a04";
		wait for Clk_period;
		Addr <=  "00100000100101";
		Trees_din <= x"ffaa20d5";
		wait for Clk_period;
		Addr <=  "00100000100110";
		Trees_din <= x"fffd20d5";
		wait for Clk_period;
		Addr <=  "00100000100111";
		Trees_din <= x"14024a08";
		wait for Clk_period;
		Addr <=  "00100000101000";
		Trees_din <= x"0e00b204";
		wait for Clk_period;
		Addr <=  "00100000101001";
		Trees_din <= x"fff720d5";
		wait for Clk_period;
		Addr <=  "00100000101010";
		Trees_din <= x"ff8b20d5";
		wait for Clk_period;
		Addr <=  "00100000101011";
		Trees_din <= x"002020d5";
		wait for Clk_period;
		Addr <=  "00100000101100";
		Trees_din <= x"08002e04";
		wait for Clk_period;
		Addr <=  "00100000101101";
		Trees_din <= x"005a20d5";
		wait for Clk_period;
		Addr <=  "00100000101110";
		Trees_din <= x"1a00c508";
		wait for Clk_period;
		Addr <=  "00100000101111";
		Trees_din <= x"17002c04";
		wait for Clk_period;
		Addr <=  "00100000110000";
		Trees_din <= x"000420d5";
		wait for Clk_period;
		Addr <=  "00100000110001";
		Trees_din <= x"ffba20d5";
		wait for Clk_period;
		Addr <=  "00100000110010";
		Trees_din <= x"0bfb2904";
		wait for Clk_period;
		Addr <=  "00100000110011";
		Trees_din <= x"fff920d5";
		wait for Clk_period;
		Addr <=  "00100000110100";
		Trees_din <= x"004920d5";
		wait for Clk_period;
		Addr <=  "00100000110101";
		Trees_din <= x"040e6444";
		wait for Clk_period;
		Addr <=  "00100000110110";
		Trees_din <= x"0afb0b20";
		wait for Clk_period;
		Addr <=  "00100000110111";
		Trees_din <= x"1200ef10";
		wait for Clk_period;
		Addr <=  "00100000111000";
		Trees_din <= x"07005808";
		wait for Clk_period;
		Addr <=  "00100000111001";
		Trees_din <= x"05fbb604";
		wait for Clk_period;
		Addr <=  "00100000111010";
		Trees_din <= x"fff12169";
		wait for Clk_period;
		Addr <=  "00100000111011";
		Trees_din <= x"ff922169";
		wait for Clk_period;
		Addr <=  "00100000111100";
		Trees_din <= x"19009904";
		wait for Clk_period;
		Addr <=  "00100000111101";
		Trees_din <= x"ffeb2169";
		wait for Clk_period;
		Addr <=  "00100000111110";
		Trees_din <= x"005e2169";
		wait for Clk_period;
		Addr <=  "00100000111111";
		Trees_din <= x"06f6f10c";
		wait for Clk_period;
		Addr <=  "00100001000000";
		Trees_din <= x"07005704";
		wait for Clk_period;
		Addr <=  "00100001000001";
		Trees_din <= x"006b2169";
		wait for Clk_period;
		Addr <=  "00100001000010";
		Trees_din <= x"13ffa204";
		wait for Clk_period;
		Addr <=  "00100001000011";
		Trees_din <= x"004c2169";
		wait for Clk_period;
		Addr <=  "00100001000100";
		Trees_din <= x"ffab2169";
		wait for Clk_period;
		Addr <=  "00100001000101";
		Trees_din <= x"ffd92169";
		wait for Clk_period;
		Addr <=  "00100001000110";
		Trees_din <= x"04fff308";
		wait for Clk_period;
		Addr <=  "00100001000111";
		Trees_din <= x"1d003b04";
		wait for Clk_period;
		Addr <=  "00100001001000";
		Trees_din <= x"ffff2169";
		wait for Clk_period;
		Addr <=  "00100001001001";
		Trees_din <= x"ff942169";
		wait for Clk_period;
		Addr <=  "00100001001010";
		Trees_din <= x"0afbee0c";
		wait for Clk_period;
		Addr <=  "00100001001011";
		Trees_din <= x"0d015004";
		wait for Clk_period;
		Addr <=  "00100001001100";
		Trees_din <= x"00012169";
		wait for Clk_period;
		Addr <=  "00100001001101";
		Trees_din <= x"10055404";
		wait for Clk_period;
		Addr <=  "00100001001110";
		Trees_din <= x"ff992169";
		wait for Clk_period;
		Addr <=  "00100001001111";
		Trees_din <= x"ffe52169";
		wait for Clk_period;
		Addr <=  "00100001010000";
		Trees_din <= x"03024708";
		wait for Clk_period;
		Addr <=  "00100001010001";
		Trees_din <= x"1c003104";
		wait for Clk_period;
		Addr <=  "00100001010010";
		Trees_din <= x"ffe62169";
		wait for Clk_period;
		Addr <=  "00100001010011";
		Trees_din <= x"00322169";
		wait for Clk_period;
		Addr <=  "00100001010100";
		Trees_din <= x"15009404";
		wait for Clk_period;
		Addr <=  "00100001010101";
		Trees_din <= x"ffbb2169";
		wait for Clk_period;
		Addr <=  "00100001010110";
		Trees_din <= x"00112169";
		wait for Clk_period;
		Addr <=  "00100001010111";
		Trees_din <= x"1a00d304";
		wait for Clk_period;
		Addr <=  "00100001011000";
		Trees_din <= x"004d2169";
		wait for Clk_period;
		Addr <=  "00100001011001";
		Trees_din <= x"00002169";
		wait for Clk_period;
		Addr <=  "00100001011010";
		Trees_din <= x"0406be2c";
		wait for Clk_period;
		Addr <=  "00100001011011";
		Trees_din <= x"0e03ab20";
		wait for Clk_period;
		Addr <=  "00100001011100";
		Trees_din <= x"06f42b04";
		wait for Clk_period;
		Addr <=  "00100001011101";
		Trees_din <= x"ff8e223d";
		wait for Clk_period;
		Addr <=  "00100001011110";
		Trees_din <= x"02ff860c";
		wait for Clk_period;
		Addr <=  "00100001011111";
		Trees_din <= x"0d03b208";
		wait for Clk_period;
		Addr <=  "00100001100000";
		Trees_din <= x"1b003604";
		wait for Clk_period;
		Addr <=  "00100001100001";
		Trees_din <= x"fffb223d";
		wait for Clk_period;
		Addr <=  "00100001100010";
		Trees_din <= x"ff85223d";
		wait for Clk_period;
		Addr <=  "00100001100011";
		Trees_din <= x"002a223d";
		wait for Clk_period;
		Addr <=  "00100001100100";
		Trees_din <= x"0afb0908";
		wait for Clk_period;
		Addr <=  "00100001100101";
		Trees_din <= x"19009b04";
		wait for Clk_period;
		Addr <=  "00100001100110";
		Trees_din <= x"ffff223d";
		wait for Clk_period;
		Addr <=  "00100001100111";
		Trees_din <= x"0060223d";
		wait for Clk_period;
		Addr <=  "00100001101000";
		Trees_din <= x"0d003404";
		wait for Clk_period;
		Addr <=  "00100001101001";
		Trees_din <= x"002c223d";
		wait for Clk_period;
		Addr <=  "00100001101010";
		Trees_din <= x"ffcd223d";
		wait for Clk_period;
		Addr <=  "00100001101011";
		Trees_din <= x"16011904";
		wait for Clk_period;
		Addr <=  "00100001101100";
		Trees_din <= x"ffd7223d";
		wait for Clk_period;
		Addr <=  "00100001101101";
		Trees_din <= x"14017704";
		wait for Clk_period;
		Addr <=  "00100001101110";
		Trees_din <= x"ffee223d";
		wait for Clk_period;
		Addr <=  "00100001101111";
		Trees_din <= x"0064223d";
		wait for Clk_period;
		Addr <=  "00100001110000";
		Trees_din <= x"16011918";
		wait for Clk_period;
		Addr <=  "00100001110001";
		Trees_din <= x"05fcab10";
		wait for Clk_period;
		Addr <=  "00100001110010";
		Trees_din <= x"05fbfd0c";
		wait for Clk_period;
		Addr <=  "00100001110011";
		Trees_din <= x"12fee404";
		wait for Clk_period;
		Addr <=  "00100001110100";
		Trees_din <= x"ffd6223d";
		wait for Clk_period;
		Addr <=  "00100001110101";
		Trees_din <= x"12020404";
		wait for Clk_period;
		Addr <=  "00100001110110";
		Trees_din <= x"0068223d";
		wait for Clk_period;
		Addr <=  "00100001110111";
		Trees_din <= x"000e223d";
		wait for Clk_period;
		Addr <=  "00100001111000";
		Trees_din <= x"ffa0223d";
		wait for Clk_period;
		Addr <=  "00100001111001";
		Trees_din <= x"09005404";
		wait for Clk_period;
		Addr <=  "00100001111010";
		Trees_din <= x"0002223d";
		wait for Clk_period;
		Addr <=  "00100001111011";
		Trees_din <= x"0073223d";
		wait for Clk_period;
		Addr <=  "00100001111100";
		Trees_din <= x"16028714";
		wait for Clk_period;
		Addr <=  "00100001111101";
		Trees_din <= x"0b04740c";
		wait for Clk_period;
		Addr <=  "00100001111110";
		Trees_din <= x"09005004";
		wait for Clk_period;
		Addr <=  "00100001111111";
		Trees_din <= x"fff5223d";
		wait for Clk_period;
		Addr <=  "00100010000000";
		Trees_din <= x"1103fb04";
		wait for Clk_period;
		Addr <=  "00100010000001";
		Trees_din <= x"ff8a223d";
		wait for Clk_period;
		Addr <=  "00100010000010";
		Trees_din <= x"ffe3223d";
		wait for Clk_period;
		Addr <=  "00100010000011";
		Trees_din <= x"0f021c04";
		wait for Clk_period;
		Addr <=  "00100010000100";
		Trees_din <= x"0041223d";
		wait for Clk_period;
		Addr <=  "00100010000101";
		Trees_din <= x"fffa223d";
		wait for Clk_period;
		Addr <=  "00100010000110";
		Trees_din <= x"030a7410";
		wait for Clk_period;
		Addr <=  "00100010000111";
		Trees_din <= x"19008c08";
		wait for Clk_period;
		Addr <=  "00100010001000";
		Trees_din <= x"15008604";
		wait for Clk_period;
		Addr <=  "00100010001001";
		Trees_din <= x"ffff223d";
		wait for Clk_period;
		Addr <=  "00100010001010";
		Trees_din <= x"0063223d";
		wait for Clk_period;
		Addr <=  "00100010001011";
		Trees_din <= x"1a00e404";
		wait for Clk_period;
		Addr <=  "00100010001100";
		Trees_din <= x"ffea223d";
		wait for Clk_period;
		Addr <=  "00100010001101";
		Trees_din <= x"0043223d";
		wait for Clk_period;
		Addr <=  "00100010001110";
		Trees_din <= x"ffc9223d";
		wait for Clk_period;
		Addr <=  "00100010001111";
		Trees_din <= x"040e643c";
		wait for Clk_period;
		Addr <=  "00100010010000";
		Trees_din <= x"07005a24";
		wait for Clk_period;
		Addr <=  "00100010010001";
		Trees_din <= x"0c03e220";
		wait for Clk_period;
		Addr <=  "00100010010010";
		Trees_din <= x"0206e310";
		wait for Clk_period;
		Addr <=  "00100010010011";
		Trees_din <= x"06f3ec08";
		wait for Clk_period;
		Addr <=  "00100010010100";
		Trees_din <= x"1e005704";
		wait for Clk_period;
		Addr <=  "00100010010101";
		Trees_din <= x"001b22c1";
		wait for Clk_period;
		Addr <=  "00100010010110";
		Trees_din <= x"ffb822c1";
		wait for Clk_period;
		Addr <=  "00100010010111";
		Trees_din <= x"1d003804";
		wait for Clk_period;
		Addr <=  "00100010011000";
		Trees_din <= x"ffc422c1";
		wait for Clk_period;
		Addr <=  "00100010011001";
		Trees_din <= x"000922c1";
		wait for Clk_period;
		Addr <=  "00100010011010";
		Trees_din <= x"1b003a08";
		wait for Clk_period;
		Addr <=  "00100010011011";
		Trees_din <= x"1b003004";
		wait for Clk_period;
		Addr <=  "00100010011100";
		Trees_din <= x"001c22c1";
		wait for Clk_period;
		Addr <=  "00100010011101";
		Trees_din <= x"ffb022c1";
		wait for Clk_period;
		Addr <=  "00100010011110";
		Trees_din <= x"1b004004";
		wait for Clk_period;
		Addr <=  "00100010011111";
		Trees_din <= x"006d22c1";
		wait for Clk_period;
		Addr <=  "00100010100000";
		Trees_din <= x"000e22c1";
		wait for Clk_period;
		Addr <=  "00100010100001";
		Trees_din <= x"004522c1";
		wait for Clk_period;
		Addr <=  "00100010100010";
		Trees_din <= x"1101260c";
		wait for Clk_period;
		Addr <=  "00100010100011";
		Trees_din <= x"13f90f04";
		wait for Clk_period;
		Addr <=  "00100010100100";
		Trees_din <= x"ffad22c1";
		wait for Clk_period;
		Addr <=  "00100010100101";
		Trees_din <= x"1a00b504";
		wait for Clk_period;
		Addr <=  "00100010100110";
		Trees_din <= x"006422c1";
		wait for Clk_period;
		Addr <=  "00100010100111";
		Trees_din <= x"000022c1";
		wait for Clk_period;
		Addr <=  "00100010101000";
		Trees_din <= x"03096508";
		wait for Clk_period;
		Addr <=  "00100010101001";
		Trees_din <= x"0d035b04";
		wait for Clk_period;
		Addr <=  "00100010101010";
		Trees_din <= x"ff9422c1";
		wait for Clk_period;
		Addr <=  "00100010101011";
		Trees_din <= x"ffe622c1";
		wait for Clk_period;
		Addr <=  "00100010101100";
		Trees_din <= x"000222c1";
		wait for Clk_period;
		Addr <=  "00100010101101";
		Trees_din <= x"1a00d304";
		wait for Clk_period;
		Addr <=  "00100010101110";
		Trees_din <= x"004822c1";
		wait for Clk_period;
		Addr <=  "00100010101111";
		Trees_din <= x"000122c1";
		wait for Clk_period;
		Addr <=  "00100010110000";
		Trees_din <= x"040a4a2c";
		wait for Clk_period;
		Addr <=  "00100010110001";
		Trees_din <= x"1a008e08";
		wait for Clk_period;
		Addr <=  "00100010110010";
		Trees_din <= x"0e00a504";
		wait for Clk_period;
		Addr <=  "00100010110011";
		Trees_din <= x"00562355";
		wait for Clk_period;
		Addr <=  "00100010110100";
		Trees_din <= x"ffd22355";
		wait for Clk_period;
		Addr <=  "00100010110101";
		Trees_din <= x"03fb1e04";
		wait for Clk_period;
		Addr <=  "00100010110110";
		Trees_din <= x"ffa22355";
		wait for Clk_period;
		Addr <=  "00100010110111";
		Trees_din <= x"1c003b10";
		wait for Clk_period;
		Addr <=  "00100010111000";
		Trees_din <= x"1b003a08";
		wait for Clk_period;
		Addr <=  "00100010111001";
		Trees_din <= x"0f004a04";
		wait for Clk_period;
		Addr <=  "00100010111010";
		Trees_din <= x"001c2355";
		wait for Clk_period;
		Addr <=  "00100010111011";
		Trees_din <= x"ffdf2355";
		wait for Clk_period;
		Addr <=  "00100010111100";
		Trees_din <= x"0e00c804";
		wait for Clk_period;
		Addr <=  "00100010111101";
		Trees_din <= x"ffe22355";
		wait for Clk_period;
		Addr <=  "00100010111110";
		Trees_din <= x"00492355";
		wait for Clk_period;
		Addr <=  "00100010111111";
		Trees_din <= x"10041408";
		wait for Clk_period;
		Addr <=  "00100011000000";
		Trees_din <= x"1a00b904";
		wait for Clk_period;
		Addr <=  "00100011000001";
		Trees_din <= x"ff8b2355";
		wait for Clk_period;
		Addr <=  "00100011000010";
		Trees_din <= x"00022355";
		wait for Clk_period;
		Addr <=  "00100011000011";
		Trees_din <= x"04077804";
		wait for Clk_period;
		Addr <=  "00100011000100";
		Trees_din <= x"ffd52355";
		wait for Clk_period;
		Addr <=  "00100011000101";
		Trees_din <= x"003c2355";
		wait for Clk_period;
		Addr <=  "00100011000110";
		Trees_din <= x"030a741c";
		wait for Clk_period;
		Addr <=  "00100011000111";
		Trees_din <= x"01068710";
		wait for Clk_period;
		Addr <=  "00100011001000";
		Trees_din <= x"07005b0c";
		wait for Clk_period;
		Addr <=  "00100011001001";
		Trees_din <= x"13004e04";
		wait for Clk_period;
		Addr <=  "00100011001010";
		Trees_din <= x"006a2355";
		wait for Clk_period;
		Addr <=  "00100011001011";
		Trees_din <= x"00fbee04";
		wait for Clk_period;
		Addr <=  "00100011001100";
		Trees_din <= x"ffd22355";
		wait for Clk_period;
		Addr <=  "00100011001101";
		Trees_din <= x"00422355";
		wait for Clk_period;
		Addr <=  "00100011001110";
		Trees_din <= x"fff32355";
		wait for Clk_period;
		Addr <=  "00100011001111";
		Trees_din <= x"13fe2d08";
		wait for Clk_period;
		Addr <=  "00100011010000";
		Trees_din <= x"13f96904";
		wait for Clk_period;
		Addr <=  "00100011010001";
		Trees_din <= x"00052355";
		wait for Clk_period;
		Addr <=  "00100011010010";
		Trees_din <= x"ffab2355";
		wait for Clk_period;
		Addr <=  "00100011010011";
		Trees_din <= x"00282355";
		wait for Clk_period;
		Addr <=  "00100011010100";
		Trees_din <= x"ffd12355";
		wait for Clk_period;
		Addr <=  "00100011010101";
		Trees_din <= x"0404aa24";
		wait for Clk_period;
		Addr <=  "00100011010110";
		Trees_din <= x"15008d10";
		wait for Clk_period;
		Addr <=  "00100011010111";
		Trees_din <= x"1c003904";
		wait for Clk_period;
		Addr <=  "00100011011000";
		Trees_din <= x"005223f9";
		wait for Clk_period;
		Addr <=  "00100011011001";
		Trees_din <= x"12019d04";
		wait for Clk_period;
		Addr <=  "00100011011010";
		Trees_din <= x"ffb023f9";
		wait for Clk_period;
		Addr <=  "00100011011011";
		Trees_din <= x"00034204";
		wait for Clk_period;
		Addr <=  "00100011011100";
		Trees_din <= x"004523f9";
		wait for Clk_period;
		Addr <=  "00100011011101";
		Trees_din <= x"ffe223f9";
		wait for Clk_period;
		Addr <=  "00100011011110";
		Trees_din <= x"15009d04";
		wait for Clk_period;
		Addr <=  "00100011011111";
		Trees_din <= x"ff9223f9";
		wait for Clk_period;
		Addr <=  "00100011100000";
		Trees_din <= x"1500a008";
		wait for Clk_period;
		Addr <=  "00100011100001";
		Trees_din <= x"07005704";
		wait for Clk_period;
		Addr <=  "00100011100010";
		Trees_din <= x"001023f9";
		wait for Clk_period;
		Addr <=  "00100011100011";
		Trees_din <= x"005223f9";
		wait for Clk_period;
		Addr <=  "00100011100100";
		Trees_din <= x"0afc5304";
		wait for Clk_period;
		Addr <=  "00100011100101";
		Trees_din <= x"fffe23f9";
		wait for Clk_period;
		Addr <=  "00100011100110";
		Trees_din <= x"ffa023f9";
		wait for Clk_period;
		Addr <=  "00100011100111";
		Trees_din <= x"0d039d24";
		wait for Clk_period;
		Addr <=  "00100011101000";
		Trees_din <= x"20040010";
		wait for Clk_period;
		Addr <=  "00100011101001";
		Trees_din <= x"1b003d0c";
		wait for Clk_period;
		Addr <=  "00100011101010";
		Trees_din <= x"1003b908";
		wait for Clk_period;
		Addr <=  "00100011101011";
		Trees_din <= x"0e008204";
		wait for Clk_period;
		Addr <=  "00100011101100";
		Trees_din <= x"001e23f9";
		wait for Clk_period;
		Addr <=  "00100011101101";
		Trees_din <= x"006123f9";
		wait for Clk_period;
		Addr <=  "00100011101110";
		Trees_din <= x"ffe423f9";
		wait for Clk_period;
		Addr <=  "00100011101111";
		Trees_din <= x"ffea23f9";
		wait for Clk_period;
		Addr <=  "00100011110000";
		Trees_din <= x"0003aa10";
		wait for Clk_period;
		Addr <=  "00100011110001";
		Trees_din <= x"06f7b308";
		wait for Clk_period;
		Addr <=  "00100011110010";
		Trees_din <= x"1d003c04";
		wait for Clk_period;
		Addr <=  "00100011110011";
		Trees_din <= x"003823f9";
		wait for Clk_period;
		Addr <=  "00100011110100";
		Trees_din <= x"fff623f9";
		wait for Clk_period;
		Addr <=  "00100011110101";
		Trees_din <= x"1c003904";
		wait for Clk_period;
		Addr <=  "00100011110110";
		Trees_din <= x"ff9b23f9";
		wait for Clk_period;
		Addr <=  "00100011110111";
		Trees_din <= x"001723f9";
		wait for Clk_period;
		Addr <=  "00100011111000";
		Trees_din <= x"ffa923f9";
		wait for Clk_period;
		Addr <=  "00100011111001";
		Trees_din <= x"09005608";
		wait for Clk_period;
		Addr <=  "00100011111010";
		Trees_din <= x"0b045804";
		wait for Clk_period;
		Addr <=  "00100011111011";
		Trees_din <= x"005723f9";
		wait for Clk_period;
		Addr <=  "00100011111100";
		Trees_din <= x"001723f9";
		wait for Clk_period;
		Addr <=  "00100011111101";
		Trees_din <= x"ffe423f9";
		wait for Clk_period;
		Addr <=  "00100011111110";
		Trees_din <= x"040e6444";
		wait for Clk_period;
		Addr <=  "00100011111111";
		Trees_din <= x"06f3d620";
		wait for Clk_period;
		Addr <=  "00100100000000";
		Trees_din <= x"02085c18";
		wait for Clk_period;
		Addr <=  "00100100000001";
		Trees_din <= x"0d028d0c";
		wait for Clk_period;
		Addr <=  "00100100000010";
		Trees_din <= x"040c1204";
		wait for Clk_period;
		Addr <=  "00100100000011";
		Trees_din <= x"ff94248d";
		wait for Clk_period;
		Addr <=  "00100100000100";
		Trees_din <= x"11015604";
		wait for Clk_period;
		Addr <=  "00100100000101";
		Trees_din <= x"ffcf248d";
		wait for Clk_period;
		Addr <=  "00100100000110";
		Trees_din <= x"0025248d";
		wait for Clk_period;
		Addr <=  "00100100000111";
		Trees_din <= x"0f003604";
		wait for Clk_period;
		Addr <=  "00100100001000";
		Trees_din <= x"ffd0248d";
		wait for Clk_period;
		Addr <=  "00100100001001";
		Trees_din <= x"10fb3704";
		wait for Clk_period;
		Addr <=  "00100100001010";
		Trees_din <= x"003f248d";
		wait for Clk_period;
		Addr <=  "00100100001011";
		Trees_din <= x"fffb248d";
		wait for Clk_period;
		Addr <=  "00100100001100";
		Trees_din <= x"1401d804";
		wait for Clk_period;
		Addr <=  "00100100001101";
		Trees_din <= x"ffe6248d";
		wait for Clk_period;
		Addr <=  "00100100001110";
		Trees_din <= x"0039248d";
		wait for Clk_period;
		Addr <=  "00100100001111";
		Trees_din <= x"09005714";
		wait for Clk_period;
		Addr <=  "00100100010000";
		Trees_din <= x"0b056f10";
		wait for Clk_period;
		Addr <=  "00100100010001";
		Trees_din <= x"1d003a08";
		wait for Clk_period;
		Addr <=  "00100100010010";
		Trees_din <= x"06f64e04";
		wait for Clk_period;
		Addr <=  "00100100010011";
		Trees_din <= x"0014248d";
		wait for Clk_period;
		Addr <=  "00100100010100";
		Trees_din <= x"ffb4248d";
		wait for Clk_period;
		Addr <=  "00100100010101";
		Trees_din <= x"07005a04";
		wait for Clk_period;
		Addr <=  "00100100010110";
		Trees_din <= x"002a248d";
		wait for Clk_period;
		Addr <=  "00100100010111";
		Trees_din <= x"ffe6248d";
		wait for Clk_period;
		Addr <=  "00100100011000";
		Trees_din <= x"ffb0248d";
		wait for Clk_period;
		Addr <=  "00100100011001";
		Trees_din <= x"0e02300c";
		wait for Clk_period;
		Addr <=  "00100100011010";
		Trees_din <= x"12028808";
		wait for Clk_period;
		Addr <=  "00100100011011";
		Trees_din <= x"0b04fc04";
		wait for Clk_period;
		Addr <=  "00100100011100";
		Trees_din <= x"ffd1248d";
		wait for Clk_period;
		Addr <=  "00100100011101";
		Trees_din <= x"002f248d";
		wait for Clk_period;
		Addr <=  "00100100011110";
		Trees_din <= x"0053248d";
		wait for Clk_period;
		Addr <=  "00100100011111";
		Trees_din <= x"ff9b248d";
		wait for Clk_period;
		Addr <=  "00100100100000";
		Trees_din <= x"05f8f704";
		wait for Clk_period;
		Addr <=  "00100100100001";
		Trees_din <= x"0000248d";
		wait for Clk_period;
		Addr <=  "00100100100010";
		Trees_din <= x"0046248d";
		wait for Clk_period;
		Addr <=  "00100100100011";
		Trees_din <= x"04065f2c";
		wait for Clk_period;
		Addr <=  "00100100100100";
		Trees_din <= x"0c024114";
		wait for Clk_period;
		Addr <=  "00100100100101";
		Trees_din <= x"09005b10";
		wait for Clk_period;
		Addr <=  "00100100100110";
		Trees_din <= x"0c004304";
		wait for Clk_period;
		Addr <=  "00100100100111";
		Trees_din <= x"000d2571";
		wait for Clk_period;
		Addr <=  "00100100101000";
		Trees_din <= x"09005408";
		wait for Clk_period;
		Addr <=  "00100100101001";
		Trees_din <= x"09005104";
		wait for Clk_period;
		Addr <=  "00100100101010";
		Trees_din <= x"ffb42571";
		wait for Clk_period;
		Addr <=  "00100100101011";
		Trees_din <= x"00132571";
		wait for Clk_period;
		Addr <=  "00100100101100";
		Trees_din <= x"ff8c2571";
		wait for Clk_period;
		Addr <=  "00100100101101";
		Trees_din <= x"00382571";
		wait for Clk_period;
		Addr <=  "00100100101110";
		Trees_din <= x"05fc1d08";
		wait for Clk_period;
		Addr <=  "00100100101111";
		Trees_din <= x"17000004";
		wait for Clk_period;
		Addr <=  "00100100110000";
		Trees_din <= x"00142571";
		wait for Clk_period;
		Addr <=  "00100100110001";
		Trees_din <= x"ffb62571";
		wait for Clk_period;
		Addr <=  "00100100110010";
		Trees_din <= x"1a00b904";
		wait for Clk_period;
		Addr <=  "00100100110011";
		Trees_din <= x"ffda2571";
		wait for Clk_period;
		Addr <=  "00100100110100";
		Trees_din <= x"0c030d08";
		wait for Clk_period;
		Addr <=  "00100100110101";
		Trees_din <= x"09005504";
		wait for Clk_period;
		Addr <=  "00100100110110";
		Trees_din <= x"001c2571";
		wait for Clk_period;
		Addr <=  "00100100110111";
		Trees_din <= x"006d2571";
		wait for Clk_period;
		Addr <=  "00100100111000";
		Trees_din <= x"00022571";
		wait for Clk_period;
		Addr <=  "00100100111001";
		Trees_din <= x"0e010920";
		wait for Clk_period;
		Addr <=  "00100100111010";
		Trees_din <= x"0e009f14";
		wait for Clk_period;
		Addr <=  "00100100111011";
		Trees_din <= x"1603e10c";
		wait for Clk_period;
		Addr <=  "00100100111100";
		Trees_din <= x"0ef97704";
		wait for Clk_period;
		Addr <=  "00100100111101";
		Trees_din <= x"ffcd2571";
		wait for Clk_period;
		Addr <=  "00100100111110";
		Trees_din <= x"0efe8604";
		wait for Clk_period;
		Addr <=  "00100100111111";
		Trees_din <= x"003d2571";
		wait for Clk_period;
		Addr <=  "00100101000000";
		Trees_din <= x"fffd2571";
		wait for Clk_period;
		Addr <=  "00100101000001";
		Trees_din <= x"00fcaf04";
		wait for Clk_period;
		Addr <=  "00100101000010";
		Trees_din <= x"00162571";
		wait for Clk_period;
		Addr <=  "00100101000011";
		Trees_din <= x"ffb32571";
		wait for Clk_period;
		Addr <=  "00100101000100";
		Trees_din <= x"0d022a08";
		wait for Clk_period;
		Addr <=  "00100101000101";
		Trees_din <= x"01056504";
		wait for Clk_period;
		Addr <=  "00100101000110";
		Trees_din <= x"00172571";
		wait for Clk_period;
		Addr <=  "00100101000111";
		Trees_din <= x"00712571";
		wait for Clk_period;
		Addr <=  "00100101001000";
		Trees_din <= x"00022571";
		wait for Clk_period;
		Addr <=  "00100101001001";
		Trees_din <= x"02ff2a10";
		wait for Clk_period;
		Addr <=  "00100101001010";
		Trees_din <= x"0f001904";
		wait for Clk_period;
		Addr <=  "00100101001011";
		Trees_din <= x"ffd32571";
		wait for Clk_period;
		Addr <=  "00100101001100";
		Trees_din <= x"1a00bf04";
		wait for Clk_period;
		Addr <=  "00100101001101";
		Trees_din <= x"ffe42571";
		wait for Clk_period;
		Addr <=  "00100101001110";
		Trees_din <= x"0d029c04";
		wait for Clk_period;
		Addr <=  "00100101001111";
		Trees_din <= x"00532571";
		wait for Clk_period;
		Addr <=  "00100101010000";
		Trees_din <= x"00122571";
		wait for Clk_period;
		Addr <=  "00100101010001";
		Trees_din <= x"01049610";
		wait for Clk_period;
		Addr <=  "00100101010010";
		Trees_din <= x"07005808";
		wait for Clk_period;
		Addr <=  "00100101010011";
		Trees_din <= x"1b003904";
		wait for Clk_period;
		Addr <=  "00100101010100";
		Trees_din <= x"ffee2571";
		wait for Clk_period;
		Addr <=  "00100101010101";
		Trees_din <= x"004d2571";
		wait for Clk_period;
		Addr <=  "00100101010110";
		Trees_din <= x"17000004";
		wait for Clk_period;
		Addr <=  "00100101010111";
		Trees_din <= x"00042571";
		wait for Clk_period;
		Addr <=  "00100101011000";
		Trees_din <= x"ffaa2571";
		wait for Clk_period;
		Addr <=  "00100101011001";
		Trees_din <= x"0c015104";
		wait for Clk_period;
		Addr <=  "00100101011010";
		Trees_din <= x"ffdb2571";
		wait for Clk_period;
		Addr <=  "00100101011011";
		Trees_din <= x"ff962571";
		wait for Clk_period;
		Addr <=  "00100101011100";
		Trees_din <= x"040e643c";
		wait for Clk_period;
		Addr <=  "00100101011101";
		Trees_din <= x"07005a28";
		wait for Clk_period;
		Addr <=  "00100101011110";
		Trees_din <= x"0bf9650c";
		wait for Clk_period;
		Addr <=  "00100101011111";
		Trees_din <= x"1e007a08";
		wait for Clk_period;
		Addr <=  "00100101100000";
		Trees_din <= x"0d01d904";
		wait for Clk_period;
		Addr <=  "00100101100001";
		Trees_din <= x"ffea25f5";
		wait for Clk_period;
		Addr <=  "00100101100010";
		Trees_din <= x"ffa225f5";
		wait for Clk_period;
		Addr <=  "00100101100011";
		Trees_din <= x"002e25f5";
		wait for Clk_period;
		Addr <=  "00100101100100";
		Trees_din <= x"1c003b10";
		wait for Clk_period;
		Addr <=  "00100101100101";
		Trees_din <= x"1b003a08";
		wait for Clk_period;
		Addr <=  "00100101100110";
		Trees_din <= x"0a02ad04";
		wait for Clk_period;
		Addr <=  "00100101100111";
		Trees_din <= x"000e25f5";
		wait for Clk_period;
		Addr <=  "00100101101000";
		Trees_din <= x"ffd025f5";
		wait for Clk_period;
		Addr <=  "00100101101001";
		Trees_din <= x"13012004";
		wait for Clk_period;
		Addr <=  "00100101101010";
		Trees_din <= x"004d25f5";
		wait for Clk_period;
		Addr <=  "00100101101011";
		Trees_din <= x"ffda25f5";
		wait for Clk_period;
		Addr <=  "00100101101100";
		Trees_din <= x"07005908";
		wait for Clk_period;
		Addr <=  "00100101101101";
		Trees_din <= x"1401f704";
		wait for Clk_period;
		Addr <=  "00100101101110";
		Trees_din <= x"fff425f5";
		wait for Clk_period;
		Addr <=  "00100101101111";
		Trees_din <= x"ffab25f5";
		wait for Clk_period;
		Addr <=  "00100101110000";
		Trees_din <= x"003a25f5";
		wait for Clk_period;
		Addr <=  "00100101110001";
		Trees_din <= x"16005e08";
		wait for Clk_period;
		Addr <=  "00100101110010";
		Trees_din <= x"1100b304";
		wait for Clk_period;
		Addr <=  "00100101110011";
		Trees_din <= x"004525f5";
		wait for Clk_period;
		Addr <=  "00100101110100";
		Trees_din <= x"ffe625f5";
		wait for Clk_period;
		Addr <=  "00100101110101";
		Trees_din <= x"0afa9a04";
		wait for Clk_period;
		Addr <=  "00100101110110";
		Trees_din <= x"001325f5";
		wait for Clk_period;
		Addr <=  "00100101110111";
		Trees_din <= x"0d035b04";
		wait for Clk_period;
		Addr <=  "00100101111000";
		Trees_din <= x"ff8b25f5";
		wait for Clk_period;
		Addr <=  "00100101111001";
		Trees_din <= x"ffe425f5";
		wait for Clk_period;
		Addr <=  "00100101111010";
		Trees_din <= x"14018004";
		wait for Clk_period;
		Addr <=  "00100101111011";
		Trees_din <= x"004825f5";
		wait for Clk_period;
		Addr <=  "00100101111100";
		Trees_din <= x"000525f5";
		wait for Clk_period;
		Addr <=  "00100101111101";
		Trees_din <= x"0404aa24";
		wait for Clk_period;
		Addr <=  "00100101111110";
		Trees_din <= x"15008d10";
		wait for Clk_period;
		Addr <=  "00100101111111";
		Trees_din <= x"1c003904";
		wait for Clk_period;
		Addr <=  "00100110000000";
		Trees_din <= x"00442691";
		wait for Clk_period;
		Addr <=  "00100110000001";
		Trees_din <= x"0d01e008";
		wait for Clk_period;
		Addr <=  "00100110000010";
		Trees_din <= x"05fe9604";
		wait for Clk_period;
		Addr <=  "00100110000011";
		Trees_din <= x"fffc2691";
		wait for Clk_period;
		Addr <=  "00100110000100";
		Trees_din <= x"00312691";
		wait for Clk_period;
		Addr <=  "00100110000101";
		Trees_din <= x"ffc22691";
		wait for Clk_period;
		Addr <=  "00100110000110";
		Trees_din <= x"15009d04";
		wait for Clk_period;
		Addr <=  "00100110000111";
		Trees_din <= x"ff992691";
		wait for Clk_period;
		Addr <=  "00100110001000";
		Trees_din <= x"1500a008";
		wait for Clk_period;
		Addr <=  "00100110001001";
		Trees_din <= x"1d004204";
		wait for Clk_period;
		Addr <=  "00100110001010";
		Trees_din <= x"000b2691";
		wait for Clk_period;
		Addr <=  "00100110001011";
		Trees_din <= x"00452691";
		wait for Clk_period;
		Addr <=  "00100110001100";
		Trees_din <= x"0afb1504";
		wait for Clk_period;
		Addr <=  "00100110001101";
		Trees_din <= x"00062691";
		wait for Clk_period;
		Addr <=  "00100110001110";
		Trees_din <= x"ffaf2691";
		wait for Clk_period;
		Addr <=  "00100110001111";
		Trees_din <= x"0d039d20";
		wait for Clk_period;
		Addr <=  "00100110010000";
		Trees_din <= x"1c002504";
		wait for Clk_period;
		Addr <=  "00100110010001";
		Trees_din <= x"ffc92691";
		wait for Clk_period;
		Addr <=  "00100110010010";
		Trees_din <= x"1c002a0c";
		wait for Clk_period;
		Addr <=  "00100110010011";
		Trees_din <= x"01fe2604";
		wait for Clk_period;
		Addr <=  "00100110010100";
		Trees_din <= x"fff52691";
		wait for Clk_period;
		Addr <=  "00100110010101";
		Trees_din <= x"04077804";
		wait for Clk_period;
		Addr <=  "00100110010110";
		Trees_din <= x"000b2691";
		wait for Clk_period;
		Addr <=  "00100110010111";
		Trees_din <= x"00622691";
		wait for Clk_period;
		Addr <=  "00100110011000";
		Trees_din <= x"00fd2508";
		wait for Clk_period;
		Addr <=  "00100110011001";
		Trees_din <= x"0c029f04";
		wait for Clk_period;
		Addr <=  "00100110011010";
		Trees_din <= x"fffb2691";
		wait for Clk_period;
		Addr <=  "00100110011011";
		Trees_din <= x"004a2691";
		wait for Clk_period;
		Addr <=  "00100110011100";
		Trees_din <= x"16000304";
		wait for Clk_period;
		Addr <=  "00100110011101";
		Trees_din <= x"00472691";
		wait for Clk_period;
		Addr <=  "00100110011110";
		Trees_din <= x"ffe02691";
		wait for Clk_period;
		Addr <=  "00100110011111";
		Trees_din <= x"09005608";
		wait for Clk_period;
		Addr <=  "00100110100000";
		Trees_din <= x"0d03c404";
		wait for Clk_period;
		Addr <=  "00100110100001";
		Trees_din <= x"00192691";
		wait for Clk_period;
		Addr <=  "00100110100010";
		Trees_din <= x"00522691";
		wait for Clk_period;
		Addr <=  "00100110100011";
		Trees_din <= x"ffe82691";
		wait for Clk_period;
		Addr <=  "00100110100100";
		Trees_din <= x"040a4a3c";
		wait for Clk_period;
		Addr <=  "00100110100101";
		Trees_din <= x"1a008e08";
		wait for Clk_period;
		Addr <=  "00100110100110";
		Trees_din <= x"15007b04";
		wait for Clk_period;
		Addr <=  "00100110100111";
		Trees_din <= x"fffb273d";
		wait for Clk_period;
		Addr <=  "00100110101000";
		Trees_din <= x"004a273d";
		wait for Clk_period;
		Addr <=  "00100110101001";
		Trees_din <= x"0d00da18";
		wait for Clk_period;
		Addr <=  "00100110101010";
		Trees_din <= x"0afac208";
		wait for Clk_period;
		Addr <=  "00100110101011";
		Trees_din <= x"1b003804";
		wait for Clk_period;
		Addr <=  "00100110101100";
		Trees_din <= x"003d273d";
		wait for Clk_period;
		Addr <=  "00100110101101";
		Trees_din <= x"0005273d";
		wait for Clk_period;
		Addr <=  "00100110101110";
		Trees_din <= x"0c008308";
		wait for Clk_period;
		Addr <=  "00100110101111";
		Trees_din <= x"1b003d04";
		wait for Clk_period;
		Addr <=  "00100110110000";
		Trees_din <= x"002a273d";
		wait for Clk_period;
		Addr <=  "00100110110001";
		Trees_din <= x"ffcb273d";
		wait for Clk_period;
		Addr <=  "00100110110010";
		Trees_din <= x"18003904";
		wait for Clk_period;
		Addr <=  "00100110110011";
		Trees_din <= x"ffe4273d";
		wait for Clk_period;
		Addr <=  "00100110110100";
		Trees_din <= x"ff93273d";
		wait for Clk_period;
		Addr <=  "00100110110101";
		Trees_din <= x"0afab10c";
		wait for Clk_period;
		Addr <=  "00100110110110";
		Trees_din <= x"1b004108";
		wait for Clk_period;
		Addr <=  "00100110110111";
		Trees_din <= x"1c002c04";
		wait for Clk_period;
		Addr <=  "00100110111000";
		Trees_din <= x"ffee273d";
		wait for Clk_period;
		Addr <=  "00100110111001";
		Trees_din <= x"ff9e273d";
		wait for Clk_period;
		Addr <=  "00100110111010";
		Trees_din <= x"0014273d";
		wait for Clk_period;
		Addr <=  "00100110111011";
		Trees_din <= x"01096908";
		wait for Clk_period;
		Addr <=  "00100110111100";
		Trees_din <= x"1900a904";
		wait for Clk_period;
		Addr <=  "00100110111101";
		Trees_din <= x"001f273d";
		wait for Clk_period;
		Addr <=  "00100110111110";
		Trees_din <= x"ffd9273d";
		wait for Clk_period;
		Addr <=  "00100110111111";
		Trees_din <= x"14012704";
		wait for Clk_period;
		Addr <=  "00100111000000";
		Trees_din <= x"ffec273d";
		wait for Clk_period;
		Addr <=  "00100111000001";
		Trees_din <= x"ffa7273d";
		wait for Clk_period;
		Addr <=  "00100111000010";
		Trees_din <= x"030a7418";
		wait for Clk_period;
		Addr <=  "00100111000011";
		Trees_din <= x"08000904";
		wait for Clk_period;
		Addr <=  "00100111000100";
		Trees_din <= x"ffe2273d";
		wait for Clk_period;
		Addr <=  "00100111000101";
		Trees_din <= x"0f003404";
		wait for Clk_period;
		Addr <=  "00100111000110";
		Trees_din <= x"ffee273d";
		wait for Clk_period;
		Addr <=  "00100111000111";
		Trees_din <= x"0f024808";
		wait for Clk_period;
		Addr <=  "00100111001000";
		Trees_din <= x"0bfa8d04";
		wait for Clk_period;
		Addr <=  "00100111001001";
		Trees_din <= x"001f273d";
		wait for Clk_period;
		Addr <=  "00100111001010";
		Trees_din <= x"006f273d";
		wait for Clk_period;
		Addr <=  "00100111001011";
		Trees_din <= x"0a028704";
		wait for Clk_period;
		Addr <=  "00100111001100";
		Trees_din <= x"0024273d";
		wait for Clk_period;
		Addr <=  "00100111001101";
		Trees_din <= x"ffd7273d";
		wait for Clk_period;
		Addr <=  "00100111001110";
		Trees_din <= x"ffd6273d";
		wait for Clk_period;
		Addr <=  "00100111001111";
		Trees_din <= x"040e643c";
		wait for Clk_period;
		Addr <=  "00100111010000";
		Trees_din <= x"07005a28";
		wait for Clk_period;
		Addr <=  "00100111010001";
		Trees_din <= x"06f4f214";
		wait for Clk_period;
		Addr <=  "00100111010010";
		Trees_din <= x"0b04820c";
		wait for Clk_period;
		Addr <=  "00100111010011";
		Trees_din <= x"02085c08";
		wait for Clk_period;
		Addr <=  "00100111010100";
		Trees_din <= x"0d039304";
		wait for Clk_period;
		Addr <=  "00100111010101";
		Trees_din <= x"ffb527c1";
		wait for Clk_period;
		Addr <=  "00100111010110";
		Trees_din <= x"003427c1";
		wait for Clk_period;
		Addr <=  "00100111010111";
		Trees_din <= x"002327c1";
		wait for Clk_period;
		Addr <=  "00100111011000";
		Trees_din <= x"02000f04";
		wait for Clk_period;
		Addr <=  "00100111011001";
		Trees_din <= x"005527c1";
		wait for Clk_period;
		Addr <=  "00100111011010";
		Trees_din <= x"fff027c1";
		wait for Clk_period;
		Addr <=  "00100111011011";
		Trees_din <= x"1a00fe10";
		wait for Clk_period;
		Addr <=  "00100111011100";
		Trees_din <= x"0afa1a08";
		wait for Clk_period;
		Addr <=  "00100111011101";
		Trees_din <= x"06f76004";
		wait for Clk_period;
		Addr <=  "00100111011110";
		Trees_din <= x"ffbf27c1";
		wait for Clk_period;
		Addr <=  "00100111011111";
		Trees_din <= x"000727c1";
		wait for Clk_period;
		Addr <=  "00100111100000";
		Trees_din <= x"06f7f304";
		wait for Clk_period;
		Addr <=  "00100111100001";
		Trees_din <= x"002527c1";
		wait for Clk_period;
		Addr <=  "00100111100010";
		Trees_din <= x"ffeb27c1";
		wait for Clk_period;
		Addr <=  "00100111100011";
		Trees_din <= x"ffc127c1";
		wait for Clk_period;
		Addr <=  "00100111100100";
		Trees_din <= x"16005e08";
		wait for Clk_period;
		Addr <=  "00100111100101";
		Trees_din <= x"1100b304";
		wait for Clk_period;
		Addr <=  "00100111100110";
		Trees_din <= x"003f27c1";
		wait for Clk_period;
		Addr <=  "00100111100111";
		Trees_din <= x"ffe827c1";
		wait for Clk_period;
		Addr <=  "00100111101000";
		Trees_din <= x"0afa9a04";
		wait for Clk_period;
		Addr <=  "00100111101001";
		Trees_din <= x"000e27c1";
		wait for Clk_period;
		Addr <=  "00100111101010";
		Trees_din <= x"0d035b04";
		wait for Clk_period;
		Addr <=  "00100111101011";
		Trees_din <= x"ff9227c1";
		wait for Clk_period;
		Addr <=  "00100111101100";
		Trees_din <= x"ffe427c1";
		wait for Clk_period;
		Addr <=  "00100111101101";
		Trees_din <= x"05f8f704";
		wait for Clk_period;
		Addr <=  "00100111101110";
		Trees_din <= x"000027c1";
		wait for Clk_period;
		Addr <=  "00100111101111";
		Trees_din <= x"004227c1";
		wait for Clk_period;
		Addr <=  "00100111110000";
		Trees_din <= x"040a4a34";
		wait for Clk_period;
		Addr <=  "00100111110001";
		Trees_din <= x"1d003604";
		wait for Clk_period;
		Addr <=  "00100111110010";
		Trees_din <= x"ffc0285d";
		wait for Clk_period;
		Addr <=  "00100111110011";
		Trees_din <= x"1c002c10";
		wait for Clk_period;
		Addr <=  "00100111110100";
		Trees_din <= x"0801fa0c";
		wait for Clk_period;
		Addr <=  "00100111110101";
		Trees_din <= x"00feb704";
		wait for Clk_period;
		Addr <=  "00100111110110";
		Trees_din <= x"fffb285d";
		wait for Clk_period;
		Addr <=  "00100111110111";
		Trees_din <= x"10047f04";
		wait for Clk_period;
		Addr <=  "00100111111000";
		Trees_din <= x"004d285d";
		wait for Clk_period;
		Addr <=  "00100111111001";
		Trees_din <= x"0005285d";
		wait for Clk_period;
		Addr <=  "00100111111010";
		Trees_din <= x"ffe4285d";
		wait for Clk_period;
		Addr <=  "00100111111011";
		Trees_din <= x"01fdd910";
		wait for Clk_period;
		Addr <=  "00100111111100";
		Trees_din <= x"14013508";
		wait for Clk_period;
		Addr <=  "00100111111101";
		Trees_din <= x"06f7b004";
		wait for Clk_period;
		Addr <=  "00100111111110";
		Trees_din <= x"ffb5285d";
		wait for Clk_period;
		Addr <=  "00100111111111";
		Trees_din <= x"0000285d";
		wait for Clk_period;
		Addr <=  "00101000000000";
		Trees_din <= x"0d018404";
		wait for Clk_period;
		Addr <=  "00101000000001";
		Trees_din <= x"ffe1285d";
		wait for Clk_period;
		Addr <=  "00101000000010";
		Trees_din <= x"005f285d";
		wait for Clk_period;
		Addr <=  "00101000000011";
		Trees_din <= x"10fbfc08";
		wait for Clk_period;
		Addr <=  "00101000000100";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00101000000101";
		Trees_din <= x"001a285d";
		wait for Clk_period;
		Addr <=  "00101000000110";
		Trees_din <= x"ffaf285d";
		wait for Clk_period;
		Addr <=  "00101000000111";
		Trees_din <= x"09005a04";
		wait for Clk_period;
		Addr <=  "00101000001000";
		Trees_din <= x"ffee285d";
		wait for Clk_period;
		Addr <=  "00101000001001";
		Trees_din <= x"0042285d";
		wait for Clk_period;
		Addr <=  "00101000001010";
		Trees_din <= x"00feb714";
		wait for Clk_period;
		Addr <=  "00101000001011";
		Trees_din <= x"0b02820c";
		wait for Clk_period;
		Addr <=  "00101000001100";
		Trees_din <= x"1e007008";
		wait for Clk_period;
		Addr <=  "00101000001101";
		Trees_din <= x"02ff2a04";
		wait for Clk_period;
		Addr <=  "00101000001110";
		Trees_din <= x"fffd285d";
		wait for Clk_period;
		Addr <=  "00101000001111";
		Trees_din <= x"ffba285d";
		wait for Clk_period;
		Addr <=  "00101000010000";
		Trees_din <= x"001e285d";
		wait for Clk_period;
		Addr <=  "00101000010001";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00101000010010";
		Trees_din <= x"004d285d";
		wait for Clk_period;
		Addr <=  "00101000010011";
		Trees_din <= x"fff7285d";
		wait for Clk_period;
		Addr <=  "00101000010100";
		Trees_din <= x"13fe8704";
		wait for Clk_period;
		Addr <=  "00101000010101";
		Trees_din <= x"000f285d";
		wait for Clk_period;
		Addr <=  "00101000010110";
		Trees_din <= x"0055285d";
		wait for Clk_period;
		Addr <=  "00101000010111";
		Trees_din <= x"0406be28";
		wait for Clk_period;
		Addr <=  "00101000011000";
		Trees_din <= x"0e03ab20";
		wait for Clk_period;
		Addr <=  "00101000011001";
		Trees_din <= x"06f42b04";
		wait for Clk_period;
		Addr <=  "00101000011010";
		Trees_din <= x"ff9f2921";
		wait for Clk_period;
		Addr <=  "00101000011011";
		Trees_din <= x"02ff860c";
		wait for Clk_period;
		Addr <=  "00101000011100";
		Trees_din <= x"1e006408";
		wait for Clk_period;
		Addr <=  "00101000011101";
		Trees_din <= x"09005504";
		wait for Clk_period;
		Addr <=  "00101000011110";
		Trees_din <= x"ffcb2921";
		wait for Clk_period;
		Addr <=  "00101000011111";
		Trees_din <= x"00362921";
		wait for Clk_period;
		Addr <=  "00101000100000";
		Trees_din <= x"ffb12921";
		wait for Clk_period;
		Addr <=  "00101000100001";
		Trees_din <= x"09005708";
		wait for Clk_period;
		Addr <=  "00101000100010";
		Trees_din <= x"03ff5404";
		wait for Clk_period;
		Addr <=  "00101000100011";
		Trees_din <= x"ffe72921";
		wait for Clk_period;
		Addr <=  "00101000100100";
		Trees_din <= x"00322921";
		wait for Clk_period;
		Addr <=  "00101000100101";
		Trees_din <= x"09005a04";
		wait for Clk_period;
		Addr <=  "00101000100110";
		Trees_din <= x"ffaa2921";
		wait for Clk_period;
		Addr <=  "00101000100111";
		Trees_din <= x"000c2921";
		wait for Clk_period;
		Addr <=  "00101000101000";
		Trees_din <= x"04045e04";
		wait for Clk_period;
		Addr <=  "00101000101001";
		Trees_din <= x"fffd2921";
		wait for Clk_period;
		Addr <=  "00101000101010";
		Trees_din <= x"003b2921";
		wait for Clk_period;
		Addr <=  "00101000101011";
		Trees_din <= x"17000014";
		wait for Clk_period;
		Addr <=  "00101000101100";
		Trees_din <= x"05f9a404";
		wait for Clk_period;
		Addr <=  "00101000101101";
		Trees_din <= x"ffea2921";
		wait for Clk_period;
		Addr <=  "00101000101110";
		Trees_din <= x"00feee08";
		wait for Clk_period;
		Addr <=  "00101000101111";
		Trees_din <= x"0307f504";
		wait for Clk_period;
		Addr <=  "00101000110000";
		Trees_din <= x"00632921";
		wait for Clk_period;
		Addr <=  "00101000110001";
		Trees_din <= x"00122921";
		wait for Clk_period;
		Addr <=  "00101000110010";
		Trees_din <= x"08017904";
		wait for Clk_period;
		Addr <=  "00101000110011";
		Trees_din <= x"ffd72921";
		wait for Clk_period;
		Addr <=  "00101000110100";
		Trees_din <= x"00312921";
		wait for Clk_period;
		Addr <=  "00101000110101";
		Trees_din <= x"16028714";
		wait for Clk_period;
		Addr <=  "00101000110110";
		Trees_din <= x"0700550c";
		wait for Clk_period;
		Addr <=  "00101000110111";
		Trees_din <= x"12024708";
		wait for Clk_period;
		Addr <=  "00101000111000";
		Trees_din <= x"14018a04";
		wait for Clk_period;
		Addr <=  "00101000111001";
		Trees_din <= x"00422921";
		wait for Clk_period;
		Addr <=  "00101000111010";
		Trees_din <= x"00082921";
		wait for Clk_period;
		Addr <=  "00101000111011";
		Trees_din <= x"ffd72921";
		wait for Clk_period;
		Addr <=  "00101000111100";
		Trees_din <= x"10fac504";
		wait for Clk_period;
		Addr <=  "00101000111101";
		Trees_din <= x"000a2921";
		wait for Clk_period;
		Addr <=  "00101000111110";
		Trees_din <= x"ff9d2921";
		wait for Clk_period;
		Addr <=  "00101000111111";
		Trees_din <= x"030a7410";
		wait for Clk_period;
		Addr <=  "00101001000000";
		Trees_din <= x"0f00ee08";
		wait for Clk_period;
		Addr <=  "00101001000001";
		Trees_din <= x"00fce804";
		wait for Clk_period;
		Addr <=  "00101001000010";
		Trees_din <= x"00302921";
		wait for Clk_period;
		Addr <=  "00101001000011";
		Trees_din <= x"ffed2921";
		wait for Clk_period;
		Addr <=  "00101001000100";
		Trees_din <= x"10fc1004";
		wait for Clk_period;
		Addr <=  "00101001000101";
		Trees_din <= x"fff42921";
		wait for Clk_period;
		Addr <=  "00101001000110";
		Trees_din <= x"00672921";
		wait for Clk_period;
		Addr <=  "00101001000111";
		Trees_din <= x"ffd92921";
		wait for Clk_period;
		Addr <=  "00101001001000";
		Trees_din <= x"0406be24";
		wait for Clk_period;
		Addr <=  "00101001001001";
		Trees_din <= x"12fe6204";
		wait for Clk_period;
		Addr <=  "00101001001010";
		Trees_din <= x"ffab29e5";
		wait for Clk_period;
		Addr <=  "00101001001011";
		Trees_din <= x"0bf95804";
		wait for Clk_period;
		Addr <=  "00101001001100";
		Trees_din <= x"ffb029e5";
		wait for Clk_period;
		Addr <=  "00101001001101";
		Trees_din <= x"0d015010";
		wait for Clk_period;
		Addr <=  "00101001001110";
		Trees_din <= x"14035d08";
		wait for Clk_period;
		Addr <=  "00101001001111";
		Trees_din <= x"03033004";
		wait for Clk_period;
		Addr <=  "00101001010000";
		Trees_din <= x"ffa129e5";
		wait for Clk_period;
		Addr <=  "00101001010001";
		Trees_din <= x"fff829e5";
		wait for Clk_period;
		Addr <=  "00101001010010";
		Trees_din <= x"1403b904";
		wait for Clk_period;
		Addr <=  "00101001010011";
		Trees_din <= x"003f29e5";
		wait for Clk_period;
		Addr <=  "00101001010100";
		Trees_din <= x"ffd929e5";
		wait for Clk_period;
		Addr <=  "00101001010101";
		Trees_din <= x"01096908";
		wait for Clk_period;
		Addr <=  "00101001010110";
		Trees_din <= x"0af83804";
		wait for Clk_period;
		Addr <=  "00101001010111";
		Trees_din <= x"ffd429e5";
		wait for Clk_period;
		Addr <=  "00101001011000";
		Trees_din <= x"003329e5";
		wait for Clk_period;
		Addr <=  "00101001011001";
		Trees_din <= x"ffcb29e5";
		wait for Clk_period;
		Addr <=  "00101001011010";
		Trees_din <= x"17000014";
		wait for Clk_period;
		Addr <=  "00101001011011";
		Trees_din <= x"0e028810";
		wait for Clk_period;
		Addr <=  "00101001011100";
		Trees_din <= x"02027c0c";
		wait for Clk_period;
		Addr <=  "00101001011101";
		Trees_din <= x"0307f508";
		wait for Clk_period;
		Addr <=  "00101001011110";
		Trees_din <= x"15008c04";
		wait for Clk_period;
		Addr <=  "00101001011111";
		Trees_din <= x"001629e5";
		wait for Clk_period;
		Addr <=  "00101001100000";
		Trees_din <= x"006229e5";
		wait for Clk_period;
		Addr <=  "00101001100001";
		Trees_din <= x"000229e5";
		wait for Clk_period;
		Addr <=  "00101001100010";
		Trees_din <= x"fff629e5";
		wait for Clk_period;
		Addr <=  "00101001100011";
		Trees_din <= x"fff429e5";
		wait for Clk_period;
		Addr <=  "00101001100100";
		Trees_din <= x"09005214";
		wait for Clk_period;
		Addr <=  "00101001100101";
		Trees_din <= x"0700580c";
		wait for Clk_period;
		Addr <=  "00101001100110";
		Trees_din <= x"09004f08";
		wait for Clk_period;
		Addr <=  "00101001100111";
		Trees_din <= x"0f006a04";
		wait for Clk_period;
		Addr <=  "00101001101000";
		Trees_din <= x"002729e5";
		wait for Clk_period;
		Addr <=  "00101001101001";
		Trees_din <= x"ffe629e5";
		wait for Clk_period;
		Addr <=  "00101001101010";
		Trees_din <= x"005229e5";
		wait for Clk_period;
		Addr <=  "00101001101011";
		Trees_din <= x"19009504";
		wait for Clk_period;
		Addr <=  "00101001101100";
		Trees_din <= x"001729e5";
		wait for Clk_period;
		Addr <=  "00101001101101";
		Trees_din <= x"ffbc29e5";
		wait for Clk_period;
		Addr <=  "00101001101110";
		Trees_din <= x"0101d10c";
		wait for Clk_period;
		Addr <=  "00101001101111";
		Trees_din <= x"09005604";
		wait for Clk_period;
		Addr <=  "00101001110000";
		Trees_din <= x"003629e5";
		wait for Clk_period;
		Addr <=  "00101001110001";
		Trees_din <= x"04086a04";
		wait for Clk_period;
		Addr <=  "00101001110010";
		Trees_din <= x"ffcc29e5";
		wait for Clk_period;
		Addr <=  "00101001110011";
		Trees_din <= x"001b29e5";
		wait for Clk_period;
		Addr <=  "00101001110100";
		Trees_din <= x"0efe8604";
		wait for Clk_period;
		Addr <=  "00101001110101";
		Trees_din <= x"002d29e5";
		wait for Clk_period;
		Addr <=  "00101001110110";
		Trees_din <= x"1500a004";
		wait for Clk_period;
		Addr <=  "00101001110111";
		Trees_din <= x"ffa829e5";
		wait for Clk_period;
		Addr <=  "00101001111000";
		Trees_din <= x"000529e5";
		wait for Clk_period;
		Addr <=  "00101001111001";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  4
        -----------
		Addr <=  "00000000000000";
		Trees_din <= x"02097678";
		wait for Clk_period;
		Addr <=  "00000000000001";
		Trees_din <= x"000ceb3c";
		wait for Clk_period;
		Addr <=  "00000000000010";
		Trees_din <= x"02050720";
		wait for Clk_period;
		Addr <=  "00000000000011";
		Trees_din <= x"02015410";
		wait for Clk_period;
		Addr <=  "00000000000100";
		Trees_din <= x"18005508";
		wait for Clk_period;
		Addr <=  "00000000000101";
		Trees_din <= x"05fc1204";
		wait for Clk_period;
		Addr <=  "00000000000110";
		Trees_din <= x"ff57016d";
		wait for Clk_period;
		Addr <=  "00000000000111";
		Trees_din <= x"ff8c016d";
		wait for Clk_period;
		Addr <=  "00000000001000";
		Trees_din <= x"0bfacb04";
		wait for Clk_period;
		Addr <=  "00000000001001";
		Trees_din <= x"0190016d";
		wait for Clk_period;
		Addr <=  "00000000001010";
		Trees_din <= x"ff71016d";
		wait for Clk_period;
		Addr <=  "00000000001011";
		Trees_din <= x"010b3208";
		wait for Clk_period;
		Addr <=  "00000000001100";
		Trees_din <= x"17008704";
		wait for Clk_period;
		Addr <=  "00000000001101";
		Trees_din <= x"ffec016d";
		wait for Clk_period;
		Addr <=  "00000000001110";
		Trees_din <= x"00d4016d";
		wait for Clk_period;
		Addr <=  "00000000001111";
		Trees_din <= x"0301f904";
		wait for Clk_period;
		Addr <=  "00000000010000";
		Trees_din <= x"ff6a016d";
		wait for Clk_period;
		Addr <=  "00000000010001";
		Trees_din <= x"00b2016d";
		wait for Clk_period;
		Addr <=  "00000000010010";
		Trees_din <= x"010db610";
		wait for Clk_period;
		Addr <=  "00000000010011";
		Trees_din <= x"02071408";
		wait for Clk_period;
		Addr <=  "00000000010100";
		Trees_din <= x"00087804";
		wait for Clk_period;
		Addr <=  "00000000010101";
		Trees_din <= x"01c1016d";
		wait for Clk_period;
		Addr <=  "00000000010110";
		Trees_din <= x"0014016d";
		wait for Clk_period;
		Addr <=  "00000000010111";
		Trees_din <= x"08036904";
		wait for Clk_period;
		Addr <=  "00000000011000";
		Trees_din <= x"02a0016d";
		wait for Clk_period;
		Addr <=  "00000000011001";
		Trees_din <= x"0000016d";
		wait for Clk_period;
		Addr <=  "00000000011010";
		Trees_din <= x"1703bc08";
		wait for Clk_period;
		Addr <=  "00000000011011";
		Trees_din <= x"05faed04";
		wait for Clk_period;
		Addr <=  "00000000011100";
		Trees_din <= x"ff78016d";
		wait for Clk_period;
		Addr <=  "00000000011101";
		Trees_din <= x"008c016d";
		wait for Clk_period;
		Addr <=  "00000000011110";
		Trees_din <= x"00c1016d";
		wait for Clk_period;
		Addr <=  "00000000011111";
		Trees_din <= x"0206e320";
		wait for Clk_period;
		Addr <=  "00000000100000";
		Trees_din <= x"03f9f210";
		wait for Clk_period;
		Addr <=  "00000000100001";
		Trees_din <= x"1f00ed08";
		wait for Clk_period;
		Addr <=  "00000000100010";
		Trees_din <= x"0a07cb04";
		wait for Clk_period;
		Addr <=  "00000000100011";
		Trees_din <= x"ff4e016d";
		wait for Clk_period;
		Addr <=  "00000000100100";
		Trees_din <= x"ffb0016d";
		wait for Clk_period;
		Addr <=  "00000000100101";
		Trees_din <= x"001be904";
		wait for Clk_period;
		Addr <=  "00000000100110";
		Trees_din <= x"0027016d";
		wait for Clk_period;
		Addr <=  "00000000100111";
		Trees_din <= x"ff8f016d";
		wait for Clk_period;
		Addr <=  "00000000101000";
		Trees_din <= x"05015d08";
		wait for Clk_period;
		Addr <=  "00000000101001";
		Trees_din <= x"0ef9b704";
		wait for Clk_period;
		Addr <=  "00000000101010";
		Trees_din <= x"ffd1016d";
		wait for Clk_period;
		Addr <=  "00000000101011";
		Trees_din <= x"ff5d016d";
		wait for Clk_period;
		Addr <=  "00000000101100";
		Trees_din <= x"1601c004";
		wait for Clk_period;
		Addr <=  "00000000101101";
		Trees_din <= x"013c016d";
		wait for Clk_period;
		Addr <=  "00000000101110";
		Trees_din <= x"ff85016d";
		wait for Clk_period;
		Addr <=  "00000000101111";
		Trees_din <= x"000f6f0c";
		wait for Clk_period;
		Addr <=  "00000000110000";
		Trees_din <= x"11ffce04";
		wait for Clk_period;
		Addr <=  "00000000110001";
		Trees_din <= x"01f8016d";
		wait for Clk_period;
		Addr <=  "00000000110010";
		Trees_din <= x"000f0704";
		wait for Clk_period;
		Addr <=  "00000000110011";
		Trees_din <= x"ff9c016d";
		wait for Clk_period;
		Addr <=  "00000000110100";
		Trees_din <= x"00b2016d";
		wait for Clk_period;
		Addr <=  "00000000110101";
		Trees_din <= x"04f95808";
		wait for Clk_period;
		Addr <=  "00000000110110";
		Trees_din <= x"20028804";
		wait for Clk_period;
		Addr <=  "00000000110111";
		Trees_din <= x"ffd0016d";
		wait for Clk_period;
		Addr <=  "00000000111000";
		Trees_din <= x"ff51016d";
		wait for Clk_period;
		Addr <=  "00000000111001";
		Trees_din <= x"03f68204";
		wait for Clk_period;
		Addr <=  "00000000111010";
		Trees_din <= x"0077016d";
		wait for Clk_period;
		Addr <=  "00000000111011";
		Trees_din <= x"ff87016d";
		wait for Clk_period;
		Addr <=  "00000000111100";
		Trees_din <= x"000e4f20";
		wait for Clk_period;
		Addr <=  "00000000111101";
		Trees_din <= x"010fa414";
		wait for Clk_period;
		Addr <=  "00000000111110";
		Trees_din <= x"020cbe10";
		wait for Clk_period;
		Addr <=  "00000000111111";
		Trees_din <= x"010b1108";
		wait for Clk_period;
		Addr <=  "00000001000000";
		Trees_din <= x"1703dc04";
		wait for Clk_period;
		Addr <=  "00000001000001";
		Trees_din <= x"0362016d";
		wait for Clk_period;
		Addr <=  "00000001000010";
		Trees_din <= x"00e2016d";
		wait for Clk_period;
		Addr <=  "00000001000011";
		Trees_din <= x"0e007604";
		wait for Clk_period;
		Addr <=  "00000001000100";
		Trees_din <= x"0016016d";
		wait for Clk_period;
		Addr <=  "00000001000101";
		Trees_din <= x"025f016d";
		wait for Clk_period;
		Addr <=  "00000001000110";
		Trees_din <= x"03fb016d";
		wait for Clk_period;
		Addr <=  "00000001000111";
		Trees_din <= x"14014e04";
		wait for Clk_period;
		Addr <=  "00000001001000";
		Trees_din <= x"ff85016d";
		wait for Clk_period;
		Addr <=  "00000001001001";
		Trees_din <= x"10ffb104";
		wait for Clk_period;
		Addr <=  "00000001001010";
		Trees_din <= x"0027016d";
		wait for Clk_period;
		Addr <=  "00000001001011";
		Trees_din <= x"0236016d";
		wait for Clk_period;
		Addr <=  "00000001001100";
		Trees_din <= x"0016761c";
		wait for Clk_period;
		Addr <=  "00000001001101";
		Trees_din <= x"020b610c";
		wait for Clk_period;
		Addr <=  "00000001001110";
		Trees_din <= x"08015b04";
		wait for Clk_period;
		Addr <=  "00000001001111";
		Trees_din <= x"ff62016d";
		wait for Clk_period;
		Addr <=  "00000001010000";
		Trees_din <= x"0c01ad04";
		wait for Clk_period;
		Addr <=  "00000001010001";
		Trees_din <= x"ff8f016d";
		wait for Clk_period;
		Addr <=  "00000001010010";
		Trees_din <= x"0164016d";
		wait for Clk_period;
		Addr <=  "00000001010011";
		Trees_din <= x"09005108";
		wait for Clk_period;
		Addr <=  "00000001010100";
		Trees_din <= x"0afccf04";
		wait for Clk_period;
		Addr <=  "00000001010101";
		Trees_din <= x"ff7a016d";
		wait for Clk_period;
		Addr <=  "00000001010110";
		Trees_din <= x"00b2016d";
		wait for Clk_period;
		Addr <=  "00000001010111";
		Trees_din <= x"0e010f04";
		wait for Clk_period;
		Addr <=  "00000001011000";
		Trees_din <= x"00f6016d";
		wait for Clk_period;
		Addr <=  "00000001011001";
		Trees_din <= x"02d1016d";
		wait for Clk_period;
		Addr <=  "00000001011010";
		Trees_din <= x"ff56016d";
		wait for Clk_period;
		Addr <=  "00000001011011";
		Trees_din <= x"02083274";
		wait for Clk_period;
		Addr <=  "00000001011100";
		Trees_din <= x"000c8c40";
		wait for Clk_period;
		Addr <=  "00000001011101";
		Trees_din <= x"0202d920";
		wait for Clk_period;
		Addr <=  "00000001011110";
		Trees_din <= x"02ff0b10";
		wait for Clk_period;
		Addr <=  "00000001011111";
		Trees_din <= x"09004008";
		wait for Clk_period;
		Addr <=  "00000001100000";
		Trees_din <= x"02fe9404";
		wait for Clk_period;
		Addr <=  "00000001100001";
		Trees_din <= x"ff8702e1";
		wait for Clk_period;
		Addr <=  "00000001100010";
		Trees_din <= x"00b002e1";
		wait for Clk_period;
		Addr <=  "00000001100011";
		Trees_din <= x"0f000004";
		wait for Clk_period;
		Addr <=  "00000001100100";
		Trees_din <= x"ffc302e1";
		wait for Clk_period;
		Addr <=  "00000001100101";
		Trees_din <= x"ff5d02e1";
		wait for Clk_period;
		Addr <=  "00000001100110";
		Trees_din <= x"05fbe008";
		wait for Clk_period;
		Addr <=  "00000001100111";
		Trees_din <= x"1d005c04";
		wait for Clk_period;
		Addr <=  "00000001101000";
		Trees_din <= x"ff8102e1";
		wait for Clk_period;
		Addr <=  "00000001101001";
		Trees_din <= x"00d502e1";
		wait for Clk_period;
		Addr <=  "00000001101010";
		Trees_din <= x"04025d04";
		wait for Clk_period;
		Addr <=  "00000001101011";
		Trees_din <= x"ff9102e1";
		wait for Clk_period;
		Addr <=  "00000001101100";
		Trees_din <= x"004e02e1";
		wait for Clk_period;
		Addr <=  "00000001101101";
		Trees_din <= x"010f7410";
		wait for Clk_period;
		Addr <=  "00000001101110";
		Trees_din <= x"02049a08";
		wait for Clk_period;
		Addr <=  "00000001101111";
		Trees_din <= x"0c030d04";
		wait for Clk_period;
		Addr <=  "00000001110000";
		Trees_din <= x"009902e1";
		wait for Clk_period;
		Addr <=  "00000001110001";
		Trees_din <= x"ff6402e1";
		wait for Clk_period;
		Addr <=  "00000001110010";
		Trees_din <= x"0801bd04";
		wait for Clk_period;
		Addr <=  "00000001110011";
		Trees_din <= x"012602e1";
		wait for Clk_period;
		Addr <=  "00000001110100";
		Trees_din <= x"006b02e1";
		wait for Clk_period;
		Addr <=  "00000001110101";
		Trees_din <= x"04022408";
		wait for Clk_period;
		Addr <=  "00000001110110";
		Trees_din <= x"1c005004";
		wait for Clk_period;
		Addr <=  "00000001110111";
		Trees_din <= x"ff6202e1";
		wait for Clk_period;
		Addr <=  "00000001111000";
		Trees_din <= x"004102e1";
		wait for Clk_period;
		Addr <=  "00000001111001";
		Trees_din <= x"0c01c804";
		wait for Clk_period;
		Addr <=  "00000001111010";
		Trees_din <= x"ffa802e1";
		wait for Clk_period;
		Addr <=  "00000001111011";
		Trees_din <= x"00ce02e1";
		wait for Clk_period;
		Addr <=  "00000001111100";
		Trees_din <= x"0014d020";
		wait for Clk_period;
		Addr <=  "00000001111101";
		Trees_din <= x"0205be10";
		wait for Clk_period;
		Addr <=  "00000001111110";
		Trees_din <= x"0501a408";
		wait for Clk_period;
		Addr <=  "00000001111111";
		Trees_din <= x"08026904";
		wait for Clk_period;
		Addr <=  "00000010000000";
		Trees_din <= x"ff5602e1";
		wait for Clk_period;
		Addr <=  "00000010000001";
		Trees_din <= x"ff9902e1";
		wait for Clk_period;
		Addr <=  "00000010000010";
		Trees_din <= x"1a00c404";
		wait for Clk_period;
		Addr <=  "00000010000011";
		Trees_din <= x"00d302e1";
		wait for Clk_period;
		Addr <=  "00000010000100";
		Trees_din <= x"ff7902e1";
		wait for Clk_period;
		Addr <=  "00000010000101";
		Trees_din <= x"13fdc608";
		wait for Clk_period;
		Addr <=  "00000010000110";
		Trees_din <= x"13f90f04";
		wait for Clk_period;
		Addr <=  "00000010000111";
		Trees_din <= x"ff7c02e1";
		wait for Clk_period;
		Addr <=  "00000010001000";
		Trees_din <= x"00a702e1";
		wait for Clk_period;
		Addr <=  "00000010001001";
		Trees_din <= x"03fae604";
		wait for Clk_period;
		Addr <=  "00000010001010";
		Trees_din <= x"ff7702e1";
		wait for Clk_period;
		Addr <=  "00000010001011";
		Trees_din <= x"002402e1";
		wait for Clk_period;
		Addr <=  "00000010001100";
		Trees_din <= x"1a01370c";
		wait for Clk_period;
		Addr <=  "00000010001101";
		Trees_din <= x"0a07cb04";
		wait for Clk_period;
		Addr <=  "00000010001110";
		Trees_din <= x"ff5502e1";
		wait for Clk_period;
		Addr <=  "00000010001111";
		Trees_din <= x"0d00a704";
		wait for Clk_period;
		Addr <=  "00000010010000";
		Trees_din <= x"004102e1";
		wait for Clk_period;
		Addr <=  "00000010010001";
		Trees_din <= x"ff8002e1";
		wait for Clk_period;
		Addr <=  "00000010010010";
		Trees_din <= x"0d013104";
		wait for Clk_period;
		Addr <=  "00000010010011";
		Trees_din <= x"004302e1";
		wait for Clk_period;
		Addr <=  "00000010010100";
		Trees_din <= x"ff9802e1";
		wait for Clk_period;
		Addr <=  "00000010010101";
		Trees_din <= x"000fd32c";
		wait for Clk_period;
		Addr <=  "00000010010110";
		Trees_din <= x"010fa41c";
		wait for Clk_period;
		Addr <=  "00000010010111";
		Trees_din <= x"000c8c0c";
		wait for Clk_period;
		Addr <=  "00000010011000";
		Trees_din <= x"11f91704";
		wait for Clk_period;
		Addr <=  "00000010011001";
		Trees_din <= x"006002e1";
		wait for Clk_period;
		Addr <=  "00000010011010";
		Trees_din <= x"0e047b04";
		wait for Clk_period;
		Addr <=  "00000010011011";
		Trees_din <= x"01a002e1";
		wait for Clk_period;
		Addr <=  "00000010011100";
		Trees_din <= x"010902e1";
		wait for Clk_period;
		Addr <=  "00000010011101";
		Trees_din <= x"03fbf608";
		wait for Clk_period;
		Addr <=  "00000010011110";
		Trees_din <= x"0107f604";
		wait for Clk_period;
		Addr <=  "00000010011111";
		Trees_din <= x"019602e1";
		wait for Clk_period;
		Addr <=  "00000010100000";
		Trees_din <= x"00a502e1";
		wait for Clk_period;
		Addr <=  "00000010100001";
		Trees_din <= x"08005104";
		wait for Clk_period;
		Addr <=  "00000010100010";
		Trees_din <= x"002602e1";
		wait for Clk_period;
		Addr <=  "00000010100011";
		Trees_din <= x"ff7602e1";
		wait for Clk_period;
		Addr <=  "00000010100100";
		Trees_din <= x"10051a0c";
		wait for Clk_period;
		Addr <=  "00000010100101";
		Trees_din <= x"18003808";
		wait for Clk_period;
		Addr <=  "00000010100110";
		Trees_din <= x"020a7304";
		wait for Clk_period;
		Addr <=  "00000010100111";
		Trees_din <= x"ffa702e1";
		wait for Clk_period;
		Addr <=  "00000010101000";
		Trees_din <= x"016102e1";
		wait for Clk_period;
		Addr <=  "00000010101001";
		Trees_din <= x"ff6b02e1";
		wait for Clk_period;
		Addr <=  "00000010101010";
		Trees_din <= x"016f02e1";
		wait for Clk_period;
		Addr <=  "00000010101011";
		Trees_din <= x"00167618";
		wait for Clk_period;
		Addr <=  "00000010101100";
		Trees_din <= x"020b610c";
		wait for Clk_period;
		Addr <=  "00000010101101";
		Trees_din <= x"1900a208";
		wait for Clk_period;
		Addr <=  "00000010101110";
		Trees_din <= x"1c004204";
		wait for Clk_period;
		Addr <=  "00000010101111";
		Trees_din <= x"ff5f02e1";
		wait for Clk_period;
		Addr <=  "00000010110000";
		Trees_din <= x"002302e1";
		wait for Clk_period;
		Addr <=  "00000010110001";
		Trees_din <= x"008f02e1";
		wait for Clk_period;
		Addr <=  "00000010110010";
		Trees_din <= x"09005104";
		wait for Clk_period;
		Addr <=  "00000010110011";
		Trees_din <= x"ff7b02e1";
		wait for Clk_period;
		Addr <=  "00000010110100";
		Trees_din <= x"06f3f704";
		wait for Clk_period;
		Addr <=  "00000010110101";
		Trees_din <= x"006302e1";
		wait for Clk_period;
		Addr <=  "00000010110110";
		Trees_din <= x"018302e1";
		wait for Clk_period;
		Addr <=  "00000010110111";
		Trees_din <= x"ff5b02e1";
		wait for Clk_period;
		Addr <=  "00000010111000";
		Trees_din <= x"02079868";
		wait for Clk_period;
		Addr <=  "00000010111001";
		Trees_din <= x"000ceb3c";
		wait for Clk_period;
		Addr <=  "00000010111010";
		Trees_din <= x"0202d920";
		wait for Clk_period;
		Addr <=  "00000010111011";
		Trees_din <= x"02ff0b10";
		wait for Clk_period;
		Addr <=  "00000010111100";
		Trees_din <= x"09004008";
		wait for Clk_period;
		Addr <=  "00000010111101";
		Trees_din <= x"02fe9404";
		wait for Clk_period;
		Addr <=  "00000010111110";
		Trees_din <= x"ff8d045d";
		wait for Clk_period;
		Addr <=  "00000010111111";
		Trees_din <= x"0099045d";
		wait for Clk_period;
		Addr <=  "00000011000000";
		Trees_din <= x"0f000004";
		wait for Clk_period;
		Addr <=  "00000011000001";
		Trees_din <= x"ffce045d";
		wait for Clk_period;
		Addr <=  "00000011000010";
		Trees_din <= x"ff63045d";
		wait for Clk_period;
		Addr <=  "00000011000011";
		Trees_din <= x"0109e308";
		wait for Clk_period;
		Addr <=  "00000011000100";
		Trees_din <= x"1c003b04";
		wait for Clk_period;
		Addr <=  "00000011000101";
		Trees_din <= x"ffb8045d";
		wait for Clk_period;
		Addr <=  "00000011000110";
		Trees_din <= x"0052045d";
		wait for Clk_period;
		Addr <=  "00000011000111";
		Trees_din <= x"03024704";
		wait for Clk_period;
		Addr <=  "00000011001000";
		Trees_din <= x"ff62045d";
		wait for Clk_period;
		Addr <=  "00000011001001";
		Trees_din <= x"003a045d";
		wait for Clk_period;
		Addr <=  "00000011001010";
		Trees_din <= x"010f7410";
		wait for Clk_period;
		Addr <=  "00000011001011";
		Trees_din <= x"0a02e908";
		wait for Clk_period;
		Addr <=  "00000011001100";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00000011001101";
		Trees_din <= x"0002045d";
		wait for Clk_period;
		Addr <=  "00000011001110";
		Trees_din <= x"0087045d";
		wait for Clk_period;
		Addr <=  "00000011001111";
		Trees_din <= x"01092404";
		wait for Clk_period;
		Addr <=  "00000011010000";
		Trees_din <= x"016c045d";
		wait for Clk_period;
		Addr <=  "00000011010001";
		Trees_din <= x"ffbe045d";
		wait for Clk_period;
		Addr <=  "00000011010010";
		Trees_din <= x"04022408";
		wait for Clk_period;
		Addr <=  "00000011010011";
		Trees_din <= x"0d038804";
		wait for Clk_period;
		Addr <=  "00000011010100";
		Trees_din <= x"ff5f045d";
		wait for Clk_period;
		Addr <=  "00000011010101";
		Trees_din <= x"ffee045d";
		wait for Clk_period;
		Addr <=  "00000011010110";
		Trees_din <= x"0060045d";
		wait for Clk_period;
		Addr <=  "00000011010111";
		Trees_din <= x"0205be18";
		wait for Clk_period;
		Addr <=  "00000011011000";
		Trees_din <= x"1f00ed10";
		wait for Clk_period;
		Addr <=  "00000011011001";
		Trees_din <= x"03f9f208";
		wait for Clk_period;
		Addr <=  "00000011011010";
		Trees_din <= x"0a07cb04";
		wait for Clk_period;
		Addr <=  "00000011011011";
		Trees_din <= x"ff59045d";
		wait for Clk_period;
		Addr <=  "00000011011100";
		Trees_din <= x"ffd2045d";
		wait for Clk_period;
		Addr <=  "00000011011101";
		Trees_din <= x"05015d04";
		wait for Clk_period;
		Addr <=  "00000011011110";
		Trees_din <= x"ff6f045d";
		wait for Clk_period;
		Addr <=  "00000011011111";
		Trees_din <= x"0063045d";
		wait for Clk_period;
		Addr <=  "00000011100000";
		Trees_din <= x"0a014804";
		wait for Clk_period;
		Addr <=  "00000011100001";
		Trees_din <= x"ffaa045d";
		wait for Clk_period;
		Addr <=  "00000011100010";
		Trees_din <= x"0044045d";
		wait for Clk_period;
		Addr <=  "00000011100011";
		Trees_din <= x"09004408";
		wait for Clk_period;
		Addr <=  "00000011100100";
		Trees_din <= x"10041904";
		wait for Clk_period;
		Addr <=  "00000011100101";
		Trees_din <= x"ffa9045d";
		wait for Clk_period;
		Addr <=  "00000011100110";
		Trees_din <= x"016b045d";
		wait for Clk_period;
		Addr <=  "00000011100111";
		Trees_din <= x"00148708";
		wait for Clk_period;
		Addr <=  "00000011101000";
		Trees_din <= x"14031604";
		wait for Clk_period;
		Addr <=  "00000011101001";
		Trees_din <= x"ff91045d";
		wait for Clk_period;
		Addr <=  "00000011101010";
		Trees_din <= x"005a045d";
		wait for Clk_period;
		Addr <=  "00000011101011";
		Trees_din <= x"ff5d045d";
		wait for Clk_period;
		Addr <=  "00000011101100";
		Trees_din <= x"000fd334";
		wait for Clk_period;
		Addr <=  "00000011101101";
		Trees_din <= x"010fa420";
		wait for Clk_period;
		Addr <=  "00000011101110";
		Trees_din <= x"020c0710";
		wait for Clk_period;
		Addr <=  "00000011101111";
		Trees_din <= x"03004908";
		wait for Clk_period;
		Addr <=  "00000011110000";
		Trees_din <= x"09005504";
		wait for Clk_period;
		Addr <=  "00000011110001";
		Trees_din <= x"0103045d";
		wait for Clk_period;
		Addr <=  "00000011110010";
		Trees_din <= x"008c045d";
		wait for Clk_period;
		Addr <=  "00000011110011";
		Trees_din <= x"19007604";
		wait for Clk_period;
		Addr <=  "00000011110100";
		Trees_din <= x"fff0045d";
		wait for Clk_period;
		Addr <=  "00000011110101";
		Trees_din <= x"014b045d";
		wait for Clk_period;
		Addr <=  "00000011110110";
		Trees_din <= x"09005d08";
		wait for Clk_period;
		Addr <=  "00000011110111";
		Trees_din <= x"0e047b04";
		wait for Clk_period;
		Addr <=  "00000011111000";
		Trees_din <= x"0131045d";
		wait for Clk_period;
		Addr <=  "00000011111001";
		Trees_din <= x"00ba045d";
		wait for Clk_period;
		Addr <=  "00000011111010";
		Trees_din <= x"00042104";
		wait for Clk_period;
		Addr <=  "00000011111011";
		Trees_din <= x"00f2045d";
		wait for Clk_period;
		Addr <=  "00000011111100";
		Trees_din <= x"ffef045d";
		wait for Clk_period;
		Addr <=  "00000011111101";
		Trees_din <= x"020a7308";
		wait for Clk_period;
		Addr <=  "00000011111110";
		Trees_din <= x"0efe8f04";
		wait for Clk_period;
		Addr <=  "00000011111111";
		Trees_din <= x"003a045d";
		wait for Clk_period;
		Addr <=  "00000100000000";
		Trees_din <= x"ff6f045d";
		wait for Clk_period;
		Addr <=  "00000100000001";
		Trees_din <= x"10028708";
		wait for Clk_period;
		Addr <=  "00000100000010";
		Trees_din <= x"15009c04";
		wait for Clk_period;
		Addr <=  "00000100000011";
		Trees_din <= x"ff96045d";
		wait for Clk_period;
		Addr <=  "00000100000100";
		Trees_din <= x"0039045d";
		wait for Clk_period;
		Addr <=  "00000100000101";
		Trees_din <= x"0143045d";
		wait for Clk_period;
		Addr <=  "00000100000110";
		Trees_din <= x"020b6114";
		wait for Clk_period;
		Addr <=  "00000100000111";
		Trees_din <= x"1c00420c";
		wait for Clk_period;
		Addr <=  "00000100001000";
		Trees_din <= x"06f94508";
		wait for Clk_period;
		Addr <=  "00000100001001";
		Trees_din <= x"1b002c04";
		wait for Clk_period;
		Addr <=  "00000100001010";
		Trees_din <= x"ffcf045d";
		wait for Clk_period;
		Addr <=  "00000100001011";
		Trees_din <= x"ff5c045d";
		wait for Clk_period;
		Addr <=  "00000100001100";
		Trees_din <= x"0024045d";
		wait for Clk_period;
		Addr <=  "00000100001101";
		Trees_din <= x"18004904";
		wait for Clk_period;
		Addr <=  "00000100001110";
		Trees_din <= x"013d045d";
		wait for Clk_period;
		Addr <=  "00000100001111";
		Trees_din <= x"ff6e045d";
		wait for Clk_period;
		Addr <=  "00000100010000";
		Trees_din <= x"0016760c";
		wait for Clk_period;
		Addr <=  "00000100010001";
		Trees_din <= x"09005104";
		wait for Clk_period;
		Addr <=  "00000100010010";
		Trees_din <= x"ff82045d";
		wait for Clk_period;
		Addr <=  "00000100010011";
		Trees_din <= x"0a00c004";
		wait for Clk_period;
		Addr <=  "00000100010100";
		Trees_din <= x"012b045d";
		wait for Clk_period;
		Addr <=  "00000100010101";
		Trees_din <= x"0039045d";
		wait for Clk_period;
		Addr <=  "00000100010110";
		Trees_din <= x"ff73045d";
		wait for Clk_period;
		Addr <=  "00000100010111";
		Trees_din <= x"02071468";
		wait for Clk_period;
		Addr <=  "00000100011000";
		Trees_din <= x"000ceb38";
		wait for Clk_period;
		Addr <=  "00000100011001";
		Trees_din <= x"02026c20";
		wait for Clk_period;
		Addr <=  "00000100011010";
		Trees_din <= x"02ff0b10";
		wait for Clk_period;
		Addr <=  "00000100011011";
		Trees_din <= x"09004008";
		wait for Clk_period;
		Addr <=  "00000100011100";
		Trees_din <= x"02fe9404";
		wait for Clk_period;
		Addr <=  "00000100011101";
		Trees_din <= x"ff9305d9";
		wait for Clk_period;
		Addr <=  "00000100011110";
		Trees_din <= x"008005d9";
		wait for Clk_period;
		Addr <=  "00000100011111";
		Trees_din <= x"0f000004";
		wait for Clk_period;
		Addr <=  "00000100100000";
		Trees_din <= x"ffda05d9";
		wait for Clk_period;
		Addr <=  "00000100100001";
		Trees_din <= x"ff6805d9";
		wait for Clk_period;
		Addr <=  "00000100100010";
		Trees_din <= x"01087508";
		wait for Clk_period;
		Addr <=  "00000100100011";
		Trees_din <= x"15009304";
		wait for Clk_period;
		Addr <=  "00000100100100";
		Trees_din <= x"003605d9";
		wait for Clk_period;
		Addr <=  "00000100100101";
		Trees_din <= x"ffab05d9";
		wait for Clk_period;
		Addr <=  "00000100100110";
		Trees_din <= x"0b04fc04";
		wait for Clk_period;
		Addr <=  "00000100100111";
		Trees_din <= x"ff5e05d9";
		wait for Clk_period;
		Addr <=  "00000100101000";
		Trees_din <= x"ffe705d9";
		wait for Clk_period;
		Addr <=  "00000100101001";
		Trees_din <= x"01107310";
		wait for Clk_period;
		Addr <=  "00000100101010";
		Trees_din <= x"08001708";
		wait for Clk_period;
		Addr <=  "00000100101011";
		Trees_din <= x"0afbee04";
		wait for Clk_period;
		Addr <=  "00000100101100";
		Trees_din <= x"004905d9";
		wait for Clk_period;
		Addr <=  "00000100101101";
		Trees_din <= x"ff7205d9";
		wait for Clk_period;
		Addr <=  "00000100101110";
		Trees_din <= x"04012004";
		wait for Clk_period;
		Addr <=  "00000100101111";
		Trees_din <= x"002d05d9";
		wait for Clk_period;
		Addr <=  "00000100110000";
		Trees_din <= x"00a405d9";
		wait for Clk_period;
		Addr <=  "00000100110001";
		Trees_din <= x"05fb5b04";
		wait for Clk_period;
		Addr <=  "00000100110010";
		Trees_din <= x"ff6305d9";
		wait for Clk_period;
		Addr <=  "00000100110011";
		Trees_din <= x"002505d9";
		wait for Clk_period;
		Addr <=  "00000100110100";
		Trees_din <= x"03f9f218";
		wait for Clk_period;
		Addr <=  "00000100110101";
		Trees_din <= x"22000110";
		wait for Clk_period;
		Addr <=  "00000100110110";
		Trees_din <= x"0a07cb08";
		wait for Clk_period;
		Addr <=  "00000100110111";
		Trees_din <= x"02067004";
		wait for Clk_period;
		Addr <=  "00000100111000";
		Trees_din <= x"ff5e05d9";
		wait for Clk_period;
		Addr <=  "00000100111001";
		Trees_din <= x"ff9805d9";
		wait for Clk_period;
		Addr <=  "00000100111010";
		Trees_din <= x"18003d04";
		wait for Clk_period;
		Addr <=  "00000100111011";
		Trees_din <= x"003e05d9";
		wait for Clk_period;
		Addr <=  "00000100111100";
		Trees_din <= x"ff9e05d9";
		wait for Clk_period;
		Addr <=  "00000100111101";
		Trees_din <= x"22000204";
		wait for Clk_period;
		Addr <=  "00000100111110";
		Trees_din <= x"009205d9";
		wait for Clk_period;
		Addr <=  "00000100111111";
		Trees_din <= x"ff7a05d9";
		wait for Clk_period;
		Addr <=  "00000101000000";
		Trees_din <= x"05015d10";
		wait for Clk_period;
		Addr <=  "00000101000001";
		Trees_din <= x"08020d08";
		wait for Clk_period;
		Addr <=  "00000101000010";
		Trees_din <= x"1500aa04";
		wait for Clk_period;
		Addr <=  "00000101000011";
		Trees_din <= x"ff5e05d9";
		wait for Clk_period;
		Addr <=  "00000101000100";
		Trees_din <= x"ffe305d9";
		wait for Clk_period;
		Addr <=  "00000101000101";
		Trees_din <= x"09005704";
		wait for Clk_period;
		Addr <=  "00000101000110";
		Trees_din <= x"ff6805d9";
		wait for Clk_period;
		Addr <=  "00000101000111";
		Trees_din <= x"00b705d9";
		wait for Clk_period;
		Addr <=  "00000101001000";
		Trees_din <= x"1601c004";
		wait for Clk_period;
		Addr <=  "00000101001001";
		Trees_din <= x"012205d9";
		wait for Clk_period;
		Addr <=  "00000101001010";
		Trees_din <= x"ff9605d9";
		wait for Clk_period;
		Addr <=  "00000101001011";
		Trees_din <= x"000fd338";
		wait for Clk_period;
		Addr <=  "00000101001100";
		Trees_din <= x"010fa420";
		wait for Clk_period;
		Addr <=  "00000101001101";
		Trees_din <= x"020c0710";
		wait for Clk_period;
		Addr <=  "00000101001110";
		Trees_din <= x"0ef94308";
		wait for Clk_period;
		Addr <=  "00000101001111";
		Trees_din <= x"03fce704";
		wait for Clk_period;
		Addr <=  "00000101010000";
		Trees_din <= x"ff4f05d9";
		wait for Clk_period;
		Addr <=  "00000101010001";
		Trees_din <= x"008805d9";
		wait for Clk_period;
		Addr <=  "00000101010010";
		Trees_din <= x"000c8c04";
		wait for Clk_period;
		Addr <=  "00000101010011";
		Trees_din <= x"00c205d9";
		wait for Clk_period;
		Addr <=  "00000101010100";
		Trees_din <= x"004d05d9";
		wait for Clk_period;
		Addr <=  "00000101010101";
		Trees_din <= x"09005d08";
		wait for Clk_period;
		Addr <=  "00000101010110";
		Trees_din <= x"0f000004";
		wait for Clk_period;
		Addr <=  "00000101010111";
		Trees_din <= x"009d05d9";
		wait for Clk_period;
		Addr <=  "00000101011000";
		Trees_din <= x"00f305d9";
		wait for Clk_period;
		Addr <=  "00000101011001";
		Trees_din <= x"00042104";
		wait for Clk_period;
		Addr <=  "00000101011010";
		Trees_din <= x"00c705d9";
		wait for Clk_period;
		Addr <=  "00000101011011";
		Trees_din <= x"ffe805d9";
		wait for Clk_period;
		Addr <=  "00000101011100";
		Trees_din <= x"020a730c";
		wait for Clk_period;
		Addr <=  "00000101011101";
		Trees_din <= x"0d038804";
		wait for Clk_period;
		Addr <=  "00000101011110";
		Trees_din <= x"ff6e05d9";
		wait for Clk_period;
		Addr <=  "00000101011111";
		Trees_din <= x"08003804";
		wait for Clk_period;
		Addr <=  "00000101100000";
		Trees_din <= x"ff9e05d9";
		wait for Clk_period;
		Addr <=  "00000101100001";
		Trees_din <= x"00c805d9";
		wait for Clk_period;
		Addr <=  "00000101100010";
		Trees_din <= x"10028708";
		wait for Clk_period;
		Addr <=  "00000101100011";
		Trees_din <= x"10f99904";
		wait for Clk_period;
		Addr <=  "00000101100100";
		Trees_din <= x"003d05d9";
		wait for Clk_period;
		Addr <=  "00000101100101";
		Trees_din <= x"ff9605d9";
		wait for Clk_period;
		Addr <=  "00000101100110";
		Trees_din <= x"010305d9";
		wait for Clk_period;
		Addr <=  "00000101100111";
		Trees_din <= x"0016761c";
		wait for Clk_period;
		Addr <=  "00000101101000";
		Trees_din <= x"020b6110";
		wait for Clk_period;
		Addr <=  "00000101101001";
		Trees_din <= x"1900a108";
		wait for Clk_period;
		Addr <=  "00000101101010";
		Trees_din <= x"0e002904";
		wait for Clk_period;
		Addr <=  "00000101101011";
		Trees_din <= x"ffed05d9";
		wait for Clk_period;
		Addr <=  "00000101101100";
		Trees_din <= x"ff6705d9";
		wait for Clk_period;
		Addr <=  "00000101101101";
		Trees_din <= x"0d01a904";
		wait for Clk_period;
		Addr <=  "00000101101110";
		Trees_din <= x"ff9805d9";
		wait for Clk_period;
		Addr <=  "00000101101111";
		Trees_din <= x"016705d9";
		wait for Clk_period;
		Addr <=  "00000101110000";
		Trees_din <= x"09005104";
		wait for Clk_period;
		Addr <=  "00000101110001";
		Trees_din <= x"ff8905d9";
		wait for Clk_period;
		Addr <=  "00000101110010";
		Trees_din <= x"12fdf604";
		wait for Clk_period;
		Addr <=  "00000101110011";
		Trees_din <= x"ff9605d9";
		wait for Clk_period;
		Addr <=  "00000101110100";
		Trees_din <= x"00bd05d9";
		wait for Clk_period;
		Addr <=  "00000101110101";
		Trees_din <= x"ff6205d9";
		wait for Clk_period;
		Addr <=  "00000101110110";
		Trees_din <= x"02068564";
		wait for Clk_period;
		Addr <=  "00000101110111";
		Trees_din <= x"000bca34";
		wait for Clk_period;
		Addr <=  "00000101111000";
		Trees_din <= x"0200e11c";
		wait for Clk_period;
		Addr <=  "00000101111001";
		Trees_din <= x"05fc120c";
		wait for Clk_period;
		Addr <=  "00000101111010";
		Trees_din <= x"1d005e08";
		wait for Clk_period;
		Addr <=  "00000101111011";
		Trees_din <= x"0f000204";
		wait for Clk_period;
		Addr <=  "00000101111100";
		Trees_din <= x"ffc9073d";
		wait for Clk_period;
		Addr <=  "00000101111101";
		Trees_din <= x"ff5e073d";
		wait for Clk_period;
		Addr <=  "00000101111110";
		Trees_din <= x"0037073d";
		wait for Clk_period;
		Addr <=  "00000101111111";
		Trees_din <= x"02fda208";
		wait for Clk_period;
		Addr <=  "00000110000000";
		Trees_din <= x"01077d04";
		wait for Clk_period;
		Addr <=  "00000110000001";
		Trees_din <= x"ff62073d";
		wait for Clk_period;
		Addr <=  "00000110000010";
		Trees_din <= x"003c073d";
		wait for Clk_period;
		Addr <=  "00000110000011";
		Trees_din <= x"04025d04";
		wait for Clk_period;
		Addr <=  "00000110000100";
		Trees_din <= x"ff79073d";
		wait for Clk_period;
		Addr <=  "00000110000101";
		Trees_din <= x"0047073d";
		wait for Clk_period;
		Addr <=  "00000110000110";
		Trees_din <= x"010ed010";
		wait for Clk_period;
		Addr <=  "00000110000111";
		Trees_din <= x"08034308";
		wait for Clk_period;
		Addr <=  "00000110001000";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00000110001001";
		Trees_din <= x"0068073d";
		wait for Clk_period;
		Addr <=  "00000110001010";
		Trees_din <= x"ffe9073d";
		wait for Clk_period;
		Addr <=  "00000110001011";
		Trees_din <= x"09004a04";
		wait for Clk_period;
		Addr <=  "00000110001100";
		Trees_din <= x"008d073d";
		wait for Clk_period;
		Addr <=  "00000110001101";
		Trees_din <= x"ff5a073d";
		wait for Clk_period;
		Addr <=  "00000110001110";
		Trees_din <= x"04022404";
		wait for Clk_period;
		Addr <=  "00000110001111";
		Trees_din <= x"ff63073d";
		wait for Clk_period;
		Addr <=  "00000110010000";
		Trees_din <= x"0058073d";
		wait for Clk_period;
		Addr <=  "00000110010001";
		Trees_din <= x"03f9f214";
		wait for Clk_period;
		Addr <=  "00000110010010";
		Trees_din <= x"1f00ed10";
		wait for Clk_period;
		Addr <=  "00000110010011";
		Trees_din <= x"02067008";
		wait for Clk_period;
		Addr <=  "00000110010100";
		Trees_din <= x"0a07cb04";
		wait for Clk_period;
		Addr <=  "00000110010101";
		Trees_din <= x"ff61073d";
		wait for Clk_period;
		Addr <=  "00000110010110";
		Trees_din <= x"ffee073d";
		wait for Clk_period;
		Addr <=  "00000110010111";
		Trees_din <= x"0c018304";
		wait for Clk_period;
		Addr <=  "00000110011000";
		Trees_din <= x"ffab073d";
		wait for Clk_period;
		Addr <=  "00000110011001";
		Trees_din <= x"0046073d";
		wait for Clk_period;
		Addr <=  "00000110011010";
		Trees_din <= x"000e073d";
		wait for Clk_period;
		Addr <=  "00000110011011";
		Trees_din <= x"02047510";
		wait for Clk_period;
		Addr <=  "00000110011100";
		Trees_din <= x"08034d08";
		wait for Clk_period;
		Addr <=  "00000110011101";
		Trees_din <= x"21000104";
		wait for Clk_period;
		Addr <=  "00000110011110";
		Trees_din <= x"ff65073d";
		wait for Clk_period;
		Addr <=  "00000110011111";
		Trees_din <= x"0055073d";
		wait for Clk_period;
		Addr <=  "00000110100000";
		Trees_din <= x"0d00f804";
		wait for Clk_period;
		Addr <=  "00000110100001";
		Trees_din <= x"ff86073d";
		wait for Clk_period;
		Addr <=  "00000110100010";
		Trees_din <= x"00f4073d";
		wait for Clk_period;
		Addr <=  "00000110100011";
		Trees_din <= x"05fb0704";
		wait for Clk_period;
		Addr <=  "00000110100100";
		Trees_din <= x"ff71073d";
		wait for Clk_period;
		Addr <=  "00000110100101";
		Trees_din <= x"0c023504";
		wait for Clk_period;
		Addr <=  "00000110100110";
		Trees_din <= x"0056073d";
		wait for Clk_period;
		Addr <=  "00000110100111";
		Trees_din <= x"01b2073d";
		wait for Clk_period;
		Addr <=  "00000110101000";
		Trees_din <= x"0011923c";
		wait for Clk_period;
		Addr <=  "00000110101001";
		Trees_din <= x"020c0720";
		wait for Clk_period;
		Addr <=  "00000110101010";
		Trees_din <= x"010f7410";
		wait for Clk_period;
		Addr <=  "00000110101011";
		Trees_din <= x"03fce708";
		wait for Clk_period;
		Addr <=  "00000110101100";
		Trees_din <= x"0ef94304";
		wait for Clk_period;
		Addr <=  "00000110101101";
		Trees_din <= x"ff5c073d";
		wait for Clk_period;
		Addr <=  "00000110101110";
		Trees_din <= x"006b073d";
		wait for Clk_period;
		Addr <=  "00000110101111";
		Trees_din <= x"01090e04";
		wait for Clk_period;
		Addr <=  "00000110110000";
		Trees_din <= x"00b4073d";
		wait for Clk_period;
		Addr <=  "00000110110001";
		Trees_din <= x"ffe0073d";
		wait for Clk_period;
		Addr <=  "00000110110010";
		Trees_din <= x"1100a908";
		wait for Clk_period;
		Addr <=  "00000110110011";
		Trees_din <= x"02089504";
		wait for Clk_period;
		Addr <=  "00000110110100";
		Trees_din <= x"ff9b073d";
		wait for Clk_period;
		Addr <=  "00000110110101";
		Trees_din <= x"00e1073d";
		wait for Clk_period;
		Addr <=  "00000110110110";
		Trees_din <= x"1a00a304";
		wait for Clk_period;
		Addr <=  "00000110110111";
		Trees_din <= x"0032073d";
		wait for Clk_period;
		Addr <=  "00000110111000";
		Trees_din <= x"ff6c073d";
		wait for Clk_period;
		Addr <=  "00000110111001";
		Trees_din <= x"07005e10";
		wait for Clk_period;
		Addr <=  "00000110111010";
		Trees_din <= x"0e047b08";
		wait for Clk_period;
		Addr <=  "00000110111011";
		Trees_din <= x"00087804";
		wait for Clk_period;
		Addr <=  "00000110111100";
		Trees_din <= x"00db073d";
		wait for Clk_period;
		Addr <=  "00000110111101";
		Trees_din <= x"00ab073d";
		wait for Clk_period;
		Addr <=  "00000110111110";
		Trees_din <= x"09004c04";
		wait for Clk_period;
		Addr <=  "00000110111111";
		Trees_din <= x"ff38073d";
		wait for Clk_period;
		Addr <=  "00000111000000";
		Trees_din <= x"00b6073d";
		wait for Clk_period;
		Addr <=  "00000111000001";
		Trees_din <= x"19008908";
		wait for Clk_period;
		Addr <=  "00000111000010";
		Trees_din <= x"03f88c04";
		wait for Clk_period;
		Addr <=  "00000111000011";
		Trees_din <= x"004f073d";
		wait for Clk_period;
		Addr <=  "00000111000100";
		Trees_din <= x"ff47073d";
		wait for Clk_period;
		Addr <=  "00000111000101";
		Trees_din <= x"00af073d";
		wait for Clk_period;
		Addr <=  "00000111000110";
		Trees_din <= x"00167610";
		wait for Clk_period;
		Addr <=  "00000111000111";
		Trees_din <= x"03f68f0c";
		wait for Clk_period;
		Addr <=  "00000111001000";
		Trees_din <= x"05f88104";
		wait for Clk_period;
		Addr <=  "00000111001001";
		Trees_din <= x"ff7a073d";
		wait for Clk_period;
		Addr <=  "00000111001010";
		Trees_din <= x"0800da04";
		wait for Clk_period;
		Addr <=  "00000111001011";
		Trees_din <= x"fff2073d";
		wait for Clk_period;
		Addr <=  "00000111001100";
		Trees_din <= x"00c6073d";
		wait for Clk_period;
		Addr <=  "00000111001101";
		Trees_din <= x"ff71073d";
		wait for Clk_period;
		Addr <=  "00000111001110";
		Trees_din <= x"ff64073d";
		wait for Clk_period;
		Addr <=  "00000111001111";
		Trees_din <= x"02068568";
		wait for Clk_period;
		Addr <=  "00000111010000";
		Trees_din <= x"000ceb3c";
		wait for Clk_period;
		Addr <=  "00000111010001";
		Trees_din <= x"02012320";
		wait for Clk_period;
		Addr <=  "00000111010010";
		Trees_din <= x"05fc1210";
		wait for Clk_period;
		Addr <=  "00000111010011";
		Trees_din <= x"1203f708";
		wait for Clk_period;
		Addr <=  "00000111010100";
		Trees_din <= x"0f000204";
		wait for Clk_period;
		Addr <=  "00000111010101";
		Trees_din <= x"ffd608b1";
		wait for Clk_period;
		Addr <=  "00000111010110";
		Trees_din <= x"ff6508b1";
		wait for Clk_period;
		Addr <=  "00000111010111";
		Trees_din <= x"0c036404";
		wait for Clk_period;
		Addr <=  "00000111011000";
		Trees_din <= x"ff8b08b1";
		wait for Clk_period;
		Addr <=  "00000111011001";
		Trees_din <= x"00c508b1";
		wait for Clk_period;
		Addr <=  "00000111011010";
		Trees_din <= x"04025d08";
		wait for Clk_period;
		Addr <=  "00000111011011";
		Trees_din <= x"04f77304";
		wait for Clk_period;
		Addr <=  "00000111011100";
		Trees_din <= x"003b08b1";
		wait for Clk_period;
		Addr <=  "00000111011101";
		Trees_din <= x"ff6108b1";
		wait for Clk_period;
		Addr <=  "00000111011110";
		Trees_din <= x"02fda204";
		wait for Clk_period;
		Addr <=  "00000111011111";
		Trees_din <= x"ff8008b1";
		wait for Clk_period;
		Addr <=  "00000111100000";
		Trees_din <= x"004008b1";
		wait for Clk_period;
		Addr <=  "00000111100001";
		Trees_din <= x"010ed010";
		wait for Clk_period;
		Addr <=  "00000111100010";
		Trees_din <= x"1d003508";
		wait for Clk_period;
		Addr <=  "00000111100011";
		Trees_din <= x"0a02f804";
		wait for Clk_period;
		Addr <=  "00000111100100";
		Trees_din <= x"00f008b1";
		wait for Clk_period;
		Addr <=  "00000111100101";
		Trees_din <= x"ff9208b1";
		wait for Clk_period;
		Addr <=  "00000111100110";
		Trees_din <= x"04f8ba04";
		wait for Clk_period;
		Addr <=  "00000111100111";
		Trees_din <= x"ff8d08b1";
		wait for Clk_period;
		Addr <=  "00000111101000";
		Trees_din <= x"002808b1";
		wait for Clk_period;
		Addr <=  "00000111101001";
		Trees_din <= x"04022408";
		wait for Clk_period;
		Addr <=  "00000111101010";
		Trees_din <= x"10f76204";
		wait for Clk_period;
		Addr <=  "00000111101011";
		Trees_din <= x"001908b1";
		wait for Clk_period;
		Addr <=  "00000111101100";
		Trees_din <= x"ff6708b1";
		wait for Clk_period;
		Addr <=  "00000111101101";
		Trees_din <= x"005c08b1";
		wait for Clk_period;
		Addr <=  "00000111101110";
		Trees_din <= x"03f9f210";
		wait for Clk_period;
		Addr <=  "00000111101111";
		Trees_din <= x"1f00ed0c";
		wait for Clk_period;
		Addr <=  "00000111110000";
		Trees_din <= x"02067008";
		wait for Clk_period;
		Addr <=  "00000111110001";
		Trees_din <= x"0a07cb04";
		wait for Clk_period;
		Addr <=  "00000111110010";
		Trees_din <= x"ff6308b1";
		wait for Clk_period;
		Addr <=  "00000111110011";
		Trees_din <= x"fffc08b1";
		wait for Clk_period;
		Addr <=  "00000111110100";
		Trees_din <= x"ffff08b1";
		wait for Clk_period;
		Addr <=  "00000111110101";
		Trees_din <= x"001708b1";
		wait for Clk_period;
		Addr <=  "00000111110110";
		Trees_din <= x"02047510";
		wait for Clk_period;
		Addr <=  "00000111110111";
		Trees_din <= x"08034d08";
		wait for Clk_period;
		Addr <=  "00000111111000";
		Trees_din <= x"1203f704";
		wait for Clk_period;
		Addr <=  "00000111111001";
		Trees_din <= x"ff6c08b1";
		wait for Clk_period;
		Addr <=  "00000111111010";
		Trees_din <= x"002008b1";
		wait for Clk_period;
		Addr <=  "00000111111011";
		Trees_din <= x"09005604";
		wait for Clk_period;
		Addr <=  "00000111111100";
		Trees_din <= x"ff9108b1";
		wait for Clk_period;
		Addr <=  "00000111111101";
		Trees_din <= x"010c08b1";
		wait for Clk_period;
		Addr <=  "00000111111110";
		Trees_din <= x"05fb0704";
		wait for Clk_period;
		Addr <=  "00000111111111";
		Trees_din <= x"ff8008b1";
		wait for Clk_period;
		Addr <=  "00001000000000";
		Trees_din <= x"04fba404";
		wait for Clk_period;
		Addr <=  "00001000000001";
		Trees_din <= x"015808b1";
		wait for Clk_period;
		Addr <=  "00001000000010";
		Trees_din <= x"000f08b1";
		wait for Clk_period;
		Addr <=  "00001000000011";
		Trees_din <= x"00119240";
		wait for Clk_period;
		Addr <=  "00001000000100";
		Trees_din <= x"020c6020";
		wait for Clk_period;
		Addr <=  "00001000000101";
		Trees_din <= x"010f7410";
		wait for Clk_period;
		Addr <=  "00001000000110";
		Trees_din <= x"17007408";
		wait for Clk_period;
		Addr <=  "00001000000111";
		Trees_din <= x"1c004d04";
		wait for Clk_period;
		Addr <=  "00001000001000";
		Trees_din <= x"009608b1";
		wait for Clk_period;
		Addr <=  "00001000001001";
		Trees_din <= x"ffc808b1";
		wait for Clk_period;
		Addr <=  "00001000001010";
		Trees_din <= x"1602c904";
		wait for Clk_period;
		Addr <=  "00001000001011";
		Trees_din <= x"ffa008b1";
		wait for Clk_period;
		Addr <=  "00001000001100";
		Trees_din <= x"006608b1";
		wait for Clk_period;
		Addr <=  "00001000001101";
		Trees_din <= x"1100a908";
		wait for Clk_period;
		Addr <=  "00001000001110";
		Trees_din <= x"02089504";
		wait for Clk_period;
		Addr <=  "00001000001111";
		Trees_din <= x"ffa308b1";
		wait for Clk_period;
		Addr <=  "00001000010000";
		Trees_din <= x"00c808b1";
		wait for Clk_period;
		Addr <=  "00001000010001";
		Trees_din <= x"0e040704";
		wait for Clk_period;
		Addr <=  "00001000010010";
		Trees_din <= x"ff6f08b1";
		wait for Clk_period;
		Addr <=  "00001000010011";
		Trees_din <= x"004108b1";
		wait for Clk_period;
		Addr <=  "00001000010100";
		Trees_din <= x"0009b110";
		wait for Clk_period;
		Addr <=  "00001000010101";
		Trees_din <= x"0e047b08";
		wait for Clk_period;
		Addr <=  "00001000010110";
		Trees_din <= x"1c005004";
		wait for Clk_period;
		Addr <=  "00001000010111";
		Trees_din <= x"00c408b1";
		wait for Clk_period;
		Addr <=  "00001000011000";
		Trees_din <= x"003008b1";
		wait for Clk_period;
		Addr <=  "00001000011001";
		Trees_din <= x"0105f904";
		wait for Clk_period;
		Addr <=  "00001000011010";
		Trees_din <= x"00b408b1";
		wait for Clk_period;
		Addr <=  "00001000011011";
		Trees_din <= x"ff7008b1";
		wait for Clk_period;
		Addr <=  "00001000011100";
		Trees_din <= x"0c025308";
		wait for Clk_period;
		Addr <=  "00001000011101";
		Trees_din <= x"0c00db04";
		wait for Clk_period;
		Addr <=  "00001000011110";
		Trees_din <= x"00b208b1";
		wait for Clk_period;
		Addr <=  "00001000011111";
		Trees_din <= x"001608b1";
		wait for Clk_period;
		Addr <=  "00001000100000";
		Trees_din <= x"0f000004";
		wait for Clk_period;
		Addr <=  "00001000100001";
		Trees_din <= x"000c08b1";
		wait for Clk_period;
		Addr <=  "00001000100010";
		Trees_din <= x"00cf08b1";
		wait for Clk_period;
		Addr <=  "00001000100011";
		Trees_din <= x"00167610";
		wait for Clk_period;
		Addr <=  "00001000100100";
		Trees_din <= x"03f68f0c";
		wait for Clk_period;
		Addr <=  "00001000100101";
		Trees_din <= x"05f88104";
		wait for Clk_period;
		Addr <=  "00001000100110";
		Trees_din <= x"ff8108b1";
		wait for Clk_period;
		Addr <=  "00001000100111";
		Trees_din <= x"0e025a04";
		wait for Clk_period;
		Addr <=  "00001000101000";
		Trees_din <= x"008408b1";
		wait for Clk_period;
		Addr <=  "00001000101001";
		Trees_din <= x"ffa808b1";
		wait for Clk_period;
		Addr <=  "00001000101010";
		Trees_din <= x"ff7708b1";
		wait for Clk_period;
		Addr <=  "00001000101011";
		Trees_din <= x"ff6808b1";
		wait for Clk_period;
		Addr <=  "00001000101100";
		Trees_din <= x"02047550";
		wait for Clk_period;
		Addr <=  "00001000101101";
		Trees_din <= x"000bca3c";
		wait for Clk_period;
		Addr <=  "00001000101110";
		Trees_din <= x"02ff0b1c";
		wait for Clk_period;
		Addr <=  "00001000101111";
		Trees_din <= x"0c031c10";
		wait for Clk_period;
		Addr <=  "00001000110000";
		Trees_din <= x"09004008";
		wait for Clk_period;
		Addr <=  "00001000110001";
		Trees_din <= x"00005104";
		wait for Clk_period;
		Addr <=  "00001000110010";
		Trees_din <= x"00800a0d";
		wait for Clk_period;
		Addr <=  "00001000110011";
		Trees_din <= x"ffa30a0d";
		wait for Clk_period;
		Addr <=  "00001000110100";
		Trees_din <= x"0f000004";
		wait for Clk_period;
		Addr <=  "00001000110101";
		Trees_din <= x"000c0a0d";
		wait for Clk_period;
		Addr <=  "00001000110110";
		Trees_din <= x"ff680a0d";
		wait for Clk_period;
		Addr <=  "00001000110111";
		Trees_din <= x"02fd5104";
		wait for Clk_period;
		Addr <=  "00001000111000";
		Trees_din <= x"ff770a0d";
		wait for Clk_period;
		Addr <=  "00001000111001";
		Trees_din <= x"02fdf604";
		wait for Clk_period;
		Addr <=  "00001000111010";
		Trees_din <= x"010d0a0d";
		wait for Clk_period;
		Addr <=  "00001000111011";
		Trees_din <= x"ff930a0d";
		wait for Clk_period;
		Addr <=  "00001000111100";
		Trees_din <= x"04012010";
		wait for Clk_period;
		Addr <=  "00001000111101";
		Trees_din <= x"04fba408";
		wait for Clk_period;
		Addr <=  "00001000111110";
		Trees_din <= x"04f8a504";
		wait for Clk_period;
		Addr <=  "00001000111111";
		Trees_din <= x"ff8c0a0d";
		wait for Clk_period;
		Addr <=  "00001001000000";
		Trees_din <= x"007d0a0d";
		wait for Clk_period;
		Addr <=  "00001001000001";
		Trees_din <= x"0e03a004";
		wait for Clk_period;
		Addr <=  "00001001000010";
		Trees_din <= x"ff7a0a0d";
		wait for Clk_period;
		Addr <=  "00001001000011";
		Trees_din <= x"003a0a0d";
		wait for Clk_period;
		Addr <=  "00001001000100";
		Trees_din <= x"0c024808";
		wait for Clk_period;
		Addr <=  "00001001000101";
		Trees_din <= x"0c01d304";
		wait for Clk_period;
		Addr <=  "00001001000110";
		Trees_din <= x"00100a0d";
		wait for Clk_period;
		Addr <=  "00001001000111";
		Trees_din <= x"00ce0a0d";
		wait for Clk_period;
		Addr <=  "00001001001000";
		Trees_din <= x"15007704";
		wait for Clk_period;
		Addr <=  "00001001001001";
		Trees_din <= x"00cf0a0d";
		wait for Clk_period;
		Addr <=  "00001001001010";
		Trees_din <= x"ffb40a0d";
		wait for Clk_period;
		Addr <=  "00001001001011";
		Trees_din <= x"1f00ed10";
		wait for Clk_period;
		Addr <=  "00001001001100";
		Trees_din <= x"03fa3604";
		wait for Clk_period;
		Addr <=  "00001001001101";
		Trees_din <= x"ff640a0d";
		wait for Clk_period;
		Addr <=  "00001001001110";
		Trees_din <= x"09005c08";
		wait for Clk_period;
		Addr <=  "00001001001111";
		Trees_din <= x"13018204";
		wait for Clk_period;
		Addr <=  "00001001010000";
		Trees_din <= x"ff6f0a0d";
		wait for Clk_period;
		Addr <=  "00001001010001";
		Trees_din <= x"00450a0d";
		wait for Clk_period;
		Addr <=  "00001001010010";
		Trees_din <= x"00a40a0d";
		wait for Clk_period;
		Addr <=  "00001001010011";
		Trees_din <= x"00270a0d";
		wait for Clk_period;
		Addr <=  "00001001010100";
		Trees_din <= x"0014ad40";
		wait for Clk_period;
		Addr <=  "00001001010101";
		Trees_din <= x"020b6120";
		wait for Clk_period;
		Addr <=  "00001001010110";
		Trees_din <= x"010f7410";
		wait for Clk_period;
		Addr <=  "00001001010111";
		Trees_din <= x"000c8c08";
		wait for Clk_period;
		Addr <=  "00001001011000";
		Trees_din <= x"0ef94304";
		wait for Clk_period;
		Addr <=  "00001001011001";
		Trees_din <= x"ff760a0d";
		wait for Clk_period;
		Addr <=  "00001001011010";
		Trees_din <= x"005f0a0d";
		wait for Clk_period;
		Addr <=  "00001001011011";
		Trees_din <= x"0efddb04";
		wait for Clk_period;
		Addr <=  "00001001011100";
		Trees_din <= x"00820a0d";
		wait for Clk_period;
		Addr <=  "00001001011101";
		Trees_din <= x"ffee0a0d";
		wait for Clk_period;
		Addr <=  "00001001011110";
		Trees_din <= x"0b028808";
		wait for Clk_period;
		Addr <=  "00001001011111";
		Trees_din <= x"1d004f04";
		wait for Clk_period;
		Addr <=  "00001001100000";
		Trees_din <= x"ff6d0a0d";
		wait for Clk_period;
		Addr <=  "00001001100001";
		Trees_din <= x"00120a0d";
		wait for Clk_period;
		Addr <=  "00001001100010";
		Trees_din <= x"05f9de04";
		wait for Clk_period;
		Addr <=  "00001001100011";
		Trees_din <= x"ffc40a0d";
		wait for Clk_period;
		Addr <=  "00001001100100";
		Trees_din <= x"00cf0a0d";
		wait for Clk_period;
		Addr <=  "00001001100101";
		Trees_din <= x"000ceb10";
		wait for Clk_period;
		Addr <=  "00001001100110";
		Trees_din <= x"06fdac08";
		wait for Clk_period;
		Addr <=  "00001001100111";
		Trees_din <= x"14000d04";
		wait for Clk_period;
		Addr <=  "00001001101000";
		Trees_din <= x"ffdc0a0d";
		wait for Clk_period;
		Addr <=  "00001001101001";
		Trees_din <= x"00a30a0d";
		wait for Clk_period;
		Addr <=  "00001001101010";
		Trees_din <= x"0d02b504";
		wait for Clk_period;
		Addr <=  "00001001101011";
		Trees_din <= x"00150a0d";
		wait for Clk_period;
		Addr <=  "00001001101100";
		Trees_din <= x"ffaf0a0d";
		wait for Clk_period;
		Addr <=  "00001001101101";
		Trees_din <= x"0c01f408";
		wait for Clk_period;
		Addr <=  "00001001101110";
		Trees_din <= x"1c002e04";
		wait for Clk_period;
		Addr <=  "00001001101111";
		Trees_din <= x"00ab0a0d";
		wait for Clk_period;
		Addr <=  "00001001110000";
		Trees_din <= x"ffda0a0d";
		wait for Clk_period;
		Addr <=  "00001001110001";
		Trees_din <= x"06f34c04";
		wait for Clk_period;
		Addr <=  "00001001110010";
		Trees_din <= x"000d0a0d";
		wait for Clk_period;
		Addr <=  "00001001110011";
		Trees_din <= x"00e40a0d";
		wait for Clk_period;
		Addr <=  "00001001110100";
		Trees_din <= x"04f81510";
		wait for Clk_period;
		Addr <=  "00001001110101";
		Trees_din <= x"020d0608";
		wait for Clk_period;
		Addr <=  "00001001110110";
		Trees_din <= x"13f83c04";
		wait for Clk_period;
		Addr <=  "00001001110111";
		Trees_din <= x"00110a0d";
		wait for Clk_period;
		Addr <=  "00001001111000";
		Trees_din <= x"ff640a0d";
		wait for Clk_period;
		Addr <=  "00001001111001";
		Trees_din <= x"18004e04";
		wait for Clk_period;
		Addr <=  "00001001111010";
		Trees_din <= x"fff10a0d";
		wait for Clk_period;
		Addr <=  "00001001111011";
		Trees_din <= x"007f0a0d";
		wait for Clk_period;
		Addr <=  "00001001111100";
		Trees_din <= x"1b003508";
		wait for Clk_period;
		Addr <=  "00001001111101";
		Trees_din <= x"06f4cb04";
		wait for Clk_period;
		Addr <=  "00001001111110";
		Trees_din <= x"00260a0d";
		wait for Clk_period;
		Addr <=  "00001001111111";
		Trees_din <= x"016f0a0d";
		wait for Clk_period;
		Addr <=  "00001010000000";
		Trees_din <= x"0101d104";
		wait for Clk_period;
		Addr <=  "00001010000001";
		Trees_din <= x"000e0a0d";
		wait for Clk_period;
		Addr <=  "00001010000010";
		Trees_din <= x"ff780a0d";
		wait for Clk_period;
		Addr <=  "00001010000011";
		Trees_din <= x"0204754c";
		wait for Clk_period;
		Addr <=  "00001010000100";
		Trees_din <= x"03fa3618";
		wait for Clk_period;
		Addr <=  "00001010000101";
		Trees_din <= x"0401a510";
		wait for Clk_period;
		Addr <=  "00001010000110";
		Trees_din <= x"1f00ed0c";
		wait for Clk_period;
		Addr <=  "00001010000111";
		Trees_din <= x"10062404";
		wait for Clk_period;
		Addr <=  "00001010001000";
		Trees_din <= x"ff630b59";
		wait for Clk_period;
		Addr <=  "00001010001001";
		Trees_din <= x"00135a04";
		wait for Clk_period;
		Addr <=  "00001010001010";
		Trees_din <= x"00490b59";
		wait for Clk_period;
		Addr <=  "00001010001011";
		Trees_din <= x"ff7a0b59";
		wait for Clk_period;
		Addr <=  "00001010001100";
		Trees_din <= x"00310b59";
		wait for Clk_period;
		Addr <=  "00001010001101";
		Trees_din <= x"1200bb04";
		wait for Clk_period;
		Addr <=  "00001010001110";
		Trees_din <= x"ffa90b59";
		wait for Clk_period;
		Addr <=  "00001010001111";
		Trees_din <= x"00d90b59";
		wait for Clk_period;
		Addr <=  "00001010010000";
		Trees_din <= x"02fe8314";
		wait for Clk_period;
		Addr <=  "00001010010001";
		Trees_din <= x"0c031c08";
		wait for Clk_period;
		Addr <=  "00001010010010";
		Trees_din <= x"0f000004";
		wait for Clk_period;
		Addr <=  "00001010010011";
		Trees_din <= x"001b0b59";
		wait for Clk_period;
		Addr <=  "00001010010100";
		Trees_din <= x"ff640b59";
		wait for Clk_period;
		Addr <=  "00001010010101";
		Trees_din <= x"02fd5104";
		wait for Clk_period;
		Addr <=  "00001010010110";
		Trees_din <= x"ff7c0b59";
		wait for Clk_period;
		Addr <=  "00001010010111";
		Trees_din <= x"0402ed04";
		wait for Clk_period;
		Addr <=  "00001010011000";
		Trees_din <= x"ffa20b59";
		wait for Clk_period;
		Addr <=  "00001010011001";
		Trees_din <= x"00f10b59";
		wait for Clk_period;
		Addr <=  "00001010011010";
		Trees_din <= x"1700f110";
		wait for Clk_period;
		Addr <=  "00001010011011";
		Trees_din <= x"08003508";
		wait for Clk_period;
		Addr <=  "00001010011100";
		Trees_din <= x"18003e04";
		wait for Clk_period;
		Addr <=  "00001010011101";
		Trees_din <= x"00ee0b59";
		wait for Clk_period;
		Addr <=  "00001010011110";
		Trees_din <= x"ffe40b59";
		wait for Clk_period;
		Addr <=  "00001010011111";
		Trees_din <= x"18005504";
		wait for Clk_period;
		Addr <=  "00001010100000";
		Trees_din <= x"ffa90b59";
		wait for Clk_period;
		Addr <=  "00001010100001";
		Trees_din <= x"00bb0b59";
		wait for Clk_period;
		Addr <=  "00001010100010";
		Trees_din <= x"17012b08";
		wait for Clk_period;
		Addr <=  "00001010100011";
		Trees_din <= x"1400db04";
		wait for Clk_period;
		Addr <=  "00001010100100";
		Trees_din <= x"ff8d0b59";
		wait for Clk_period;
		Addr <=  "00001010100101";
		Trees_din <= x"01af0b59";
		wait for Clk_period;
		Addr <=  "00001010100110";
		Trees_din <= x"00fae404";
		wait for Clk_period;
		Addr <=  "00001010100111";
		Trees_din <= x"00be0b59";
		wait for Clk_period;
		Addr <=  "00001010101000";
		Trees_din <= x"ffe70b59";
		wait for Clk_period;
		Addr <=  "00001010101001";
		Trees_din <= x"0014ad3c";
		wait for Clk_period;
		Addr <=  "00001010101010";
		Trees_din <= x"020b6120";
		wait for Clk_period;
		Addr <=  "00001010101011";
		Trees_din <= x"0104ee10";
		wait for Clk_period;
		Addr <=  "00001010101100";
		Trees_din <= x"16015608";
		wait for Clk_period;
		Addr <=  "00001010101101";
		Trees_din <= x"13ffca04";
		wait for Clk_period;
		Addr <=  "00001010101110";
		Trees_din <= x"00d80b59";
		wait for Clk_period;
		Addr <=  "00001010101111";
		Trees_din <= x"fffb0b59";
		wait for Clk_period;
		Addr <=  "00001010110000";
		Trees_din <= x"10020304";
		wait for Clk_period;
		Addr <=  "00001010110001";
		Trees_din <= x"00810b59";
		wait for Clk_period;
		Addr <=  "00001010110010";
		Trees_din <= x"00080b59";
		wait for Clk_period;
		Addr <=  "00001010110011";
		Trees_din <= x"0f036f08";
		wait for Clk_period;
		Addr <=  "00001010110100";
		Trees_din <= x"0f02ce04";
		wait for Clk_period;
		Addr <=  "00001010110101";
		Trees_din <= x"00190b59";
		wait for Clk_period;
		Addr <=  "00001010110110";
		Trees_din <= x"00ca0b59";
		wait for Clk_period;
		Addr <=  "00001010110111";
		Trees_din <= x"1c002e04";
		wait for Clk_period;
		Addr <=  "00001010111000";
		Trees_din <= x"00da0b59";
		wait for Clk_period;
		Addr <=  "00001010111001";
		Trees_din <= x"ff880b59";
		wait for Clk_period;
		Addr <=  "00001010111010";
		Trees_din <= x"0211fd10";
		wait for Clk_period;
		Addr <=  "00001010111011";
		Trees_din <= x"1102a908";
		wait for Clk_period;
		Addr <=  "00001010111100";
		Trees_din <= x"06fdac04";
		wait for Clk_period;
		Addr <=  "00001010111101";
		Trees_din <= x"00850b59";
		wait for Clk_period;
		Addr <=  "00001010111110";
		Trees_din <= x"ff980b59";
		wait for Clk_period;
		Addr <=  "00001010111111";
		Trees_din <= x"11033e04";
		wait for Clk_period;
		Addr <=  "00001011000000";
		Trees_din <= x"ffcb0b59";
		wait for Clk_period;
		Addr <=  "00001011000001";
		Trees_din <= x"00790b59";
		wait for Clk_period;
		Addr <=  "00001011000010";
		Trees_din <= x"19007404";
		wait for Clk_period;
		Addr <=  "00001011000011";
		Trees_din <= x"ffcd0b59";
		wait for Clk_period;
		Addr <=  "00001011000100";
		Trees_din <= x"000fd304";
		wait for Clk_period;
		Addr <=  "00001011000101";
		Trees_din <= x"00b60b59";
		wait for Clk_period;
		Addr <=  "00001011000110";
		Trees_din <= x"fffb0b59";
		wait for Clk_period;
		Addr <=  "00001011000111";
		Trees_din <= x"04f81510";
		wait for Clk_period;
		Addr <=  "00001011001000";
		Trees_din <= x"020d0608";
		wait for Clk_period;
		Addr <=  "00001011001001";
		Trees_din <= x"12fd0d04";
		wait for Clk_period;
		Addr <=  "00001011001010";
		Trees_din <= x"001e0b59";
		wait for Clk_period;
		Addr <=  "00001011001011";
		Trees_din <= x"ff670b59";
		wait for Clk_period;
		Addr <=  "00001011001100";
		Trees_din <= x"0bf95804";
		wait for Clk_period;
		Addr <=  "00001011001101";
		Trees_din <= x"00730b59";
		wait for Clk_period;
		Addr <=  "00001011001110";
		Trees_din <= x"fff70b59";
		wait for Clk_period;
		Addr <=  "00001011001111";
		Trees_din <= x"1b003508";
		wait for Clk_period;
		Addr <=  "00001011010000";
		Trees_din <= x"0bfa8104";
		wait for Clk_period;
		Addr <=  "00001011010001";
		Trees_din <= x"015a0b59";
		wait for Clk_period;
		Addr <=  "00001011010010";
		Trees_din <= x"001e0b59";
		wait for Clk_period;
		Addr <=  "00001011010011";
		Trees_din <= x"17018e04";
		wait for Clk_period;
		Addr <=  "00001011010100";
		Trees_din <= x"ff800b59";
		wait for Clk_period;
		Addr <=  "00001011010101";
		Trees_din <= x"000d0b59";
		wait for Clk_period;
		Addr <=  "00001011010110";
		Trees_din <= x"0204754c";
		wait for Clk_period;
		Addr <=  "00001011010111";
		Trees_din <= x"03fa3618";
		wait for Clk_period;
		Addr <=  "00001011011000";
		Trees_din <= x"0401a510";
		wait for Clk_period;
		Addr <=  "00001011011001";
		Trees_din <= x"1f00ed0c";
		wait for Clk_period;
		Addr <=  "00001011011010";
		Trees_din <= x"10062404";
		wait for Clk_period;
		Addr <=  "00001011011011";
		Trees_din <= x"ff640c6d";
		wait for Clk_period;
		Addr <=  "00001011011100";
		Trees_din <= x"02fe4f04";
		wait for Clk_period;
		Addr <=  "00001011011101";
		Trees_din <= x"00480c6d";
		wait for Clk_period;
		Addr <=  "00001011011110";
		Trees_din <= x"ff800c6d";
		wait for Clk_period;
		Addr <=  "00001011011111";
		Trees_din <= x"00370c6d";
		wait for Clk_period;
		Addr <=  "00001011100000";
		Trees_din <= x"0d012804";
		wait for Clk_period;
		Addr <=  "00001011100001";
		Trees_din <= x"ffa80c6d";
		wait for Clk_period;
		Addr <=  "00001011100010";
		Trees_din <= x"00d70c6d";
		wait for Clk_period;
		Addr <=  "00001011100011";
		Trees_din <= x"02fe8314";
		wait for Clk_period;
		Addr <=  "00001011100100";
		Trees_din <= x"0c031c08";
		wait for Clk_period;
		Addr <=  "00001011100101";
		Trees_din <= x"0f000004";
		wait for Clk_period;
		Addr <=  "00001011100110";
		Trees_din <= x"001f0c6d";
		wait for Clk_period;
		Addr <=  "00001011100111";
		Trees_din <= x"ff660c6d";
		wait for Clk_period;
		Addr <=  "00001011101000";
		Trees_din <= x"02fd5104";
		wait for Clk_period;
		Addr <=  "00001011101001";
		Trees_din <= x"ff810c6d";
		wait for Clk_period;
		Addr <=  "00001011101010";
		Trees_din <= x"12012804";
		wait for Clk_period;
		Addr <=  "00001011101011";
		Trees_din <= x"00d40c6d";
		wait for Clk_period;
		Addr <=  "00001011101100";
		Trees_din <= x"ffa00c6d";
		wait for Clk_period;
		Addr <=  "00001011101101";
		Trees_din <= x"1700f110";
		wait for Clk_period;
		Addr <=  "00001011101110";
		Trees_din <= x"04022408";
		wait for Clk_period;
		Addr <=  "00001011101111";
		Trees_din <= x"0803b604";
		wait for Clk_period;
		Addr <=  "00001011110000";
		Trees_din <= x"ff960c6d";
		wait for Clk_period;
		Addr <=  "00001011110001";
		Trees_din <= x"00860c6d";
		wait for Clk_period;
		Addr <=  "00001011110010";
		Trees_din <= x"14015104";
		wait for Clk_period;
		Addr <=  "00001011110011";
		Trees_din <= x"ff660c6d";
		wait for Clk_period;
		Addr <=  "00001011110100";
		Trees_din <= x"00250c6d";
		wait for Clk_period;
		Addr <=  "00001011110101";
		Trees_din <= x"0e045008";
		wait for Clk_period;
		Addr <=  "00001011110110";
		Trees_din <= x"17011204";
		wait for Clk_period;
		Addr <=  "00001011110111";
		Trees_din <= x"00d70c6d";
		wait for Clk_period;
		Addr <=  "00001011111000";
		Trees_din <= x"fff40c6d";
		wait for Clk_period;
		Addr <=  "00001011111001";
		Trees_din <= x"18003c04";
		wait for Clk_period;
		Addr <=  "00001011111010";
		Trees_din <= x"00070c6d";
		wait for Clk_period;
		Addr <=  "00001011111011";
		Trees_din <= x"01bf0c6d";
		wait for Clk_period;
		Addr <=  "00001011111100";
		Trees_din <= x"00167634";
		wait for Clk_period;
		Addr <=  "00001011111101";
		Trees_din <= x"020e1a20";
		wait for Clk_period;
		Addr <=  "00001011111110";
		Trees_din <= x"0e024610";
		wait for Clk_period;
		Addr <=  "00001011111111";
		Trees_din <= x"1102c608";
		wait for Clk_period;
		Addr <=  "00001100000000";
		Trees_din <= x"000ceb04";
		wait for Clk_period;
		Addr <=  "00001100000001";
		Trees_din <= x"004e0c6d";
		wait for Clk_period;
		Addr <=  "00001100000010";
		Trees_din <= x"000b0c6d";
		wait for Clk_period;
		Addr <=  "00001100000011";
		Trees_din <= x"010c6804";
		wait for Clk_period;
		Addr <=  "00001100000100";
		Trees_din <= x"00e50c6d";
		wait for Clk_period;
		Addr <=  "00001100000101";
		Trees_din <= x"ffc90c6d";
		wait for Clk_period;
		Addr <=  "00001100000110";
		Trees_din <= x"06f73b08";
		wait for Clk_period;
		Addr <=  "00001100000111";
		Trees_din <= x"010bb604";
		wait for Clk_period;
		Addr <=  "00001100001000";
		Trees_din <= x"00120c6d";
		wait for Clk_period;
		Addr <=  "00001100001001";
		Trees_din <= x"ff7d0c6d";
		wait for Clk_period;
		Addr <=  "00001100001010";
		Trees_din <= x"05f6de04";
		wait for Clk_period;
		Addr <=  "00001100001011";
		Trees_din <= x"ff7c0c6d";
		wait for Clk_period;
		Addr <=  "00001100001100";
		Trees_din <= x"00890c6d";
		wait for Clk_period;
		Addr <=  "00001100001101";
		Trees_din <= x"010f740c";
		wait for Clk_period;
		Addr <=  "00001100001110";
		Trees_din <= x"09005d08";
		wait for Clk_period;
		Addr <=  "00001100001111";
		Trees_din <= x"0e06a204";
		wait for Clk_period;
		Addr <=  "00001100010000";
		Trees_din <= x"00960c6d";
		wait for Clk_period;
		Addr <=  "00001100010001";
		Trees_din <= x"ffe10c6d";
		wait for Clk_period;
		Addr <=  "00001100010010";
		Trees_din <= x"ffdc0c6d";
		wait for Clk_period;
		Addr <=  "00001100010011";
		Trees_din <= x"0f000104";
		wait for Clk_period;
		Addr <=  "00001100010100";
		Trees_din <= x"00420c6d";
		wait for Clk_period;
		Addr <=  "00001100010101";
		Trees_din <= x"ff800c6d";
		wait for Clk_period;
		Addr <=  "00001100010110";
		Trees_din <= x"04f81504";
		wait for Clk_period;
		Addr <=  "00001100010111";
		Trees_din <= x"ff6c0c6d";
		wait for Clk_period;
		Addr <=  "00001100011000";
		Trees_din <= x"16017504";
		wait for Clk_period;
		Addr <=  "00001100011001";
		Trees_din <= x"00da0c6d";
		wait for Clk_period;
		Addr <=  "00001100011010";
		Trees_din <= x"ffab0c6d";
		wait for Clk_period;
		Addr <=  "00001100011011";
		Trees_din <= x"02047554";
		wait for Clk_period;
		Addr <=  "00001100011100";
		Trees_din <= x"03fa3618";
		wait for Clk_period;
		Addr <=  "00001100011101";
		Trees_din <= x"0401a510";
		wait for Clk_period;
		Addr <=  "00001100011110";
		Trees_din <= x"1f00ed0c";
		wait for Clk_period;
		Addr <=  "00001100011111";
		Trees_din <= x"10062404";
		wait for Clk_period;
		Addr <=  "00001100100000";
		Trees_din <= x"ff650d89";
		wait for Clk_period;
		Addr <=  "00001100100001";
		Trees_din <= x"0c02ae04";
		wait for Clk_period;
		Addr <=  "00001100100010";
		Trees_din <= x"ff870d89";
		wait for Clk_period;
		Addr <=  "00001100100011";
		Trees_din <= x"00460d89";
		wait for Clk_period;
		Addr <=  "00001100100100";
		Trees_din <= x"003e0d89";
		wait for Clk_period;
		Addr <=  "00001100100101";
		Trees_din <= x"13fe9b04";
		wait for Clk_period;
		Addr <=  "00001100100110";
		Trees_din <= x"ffa90d89";
		wait for Clk_period;
		Addr <=  "00001100100111";
		Trees_din <= x"00d10d89";
		wait for Clk_period;
		Addr <=  "00001100101000";
		Trees_din <= x"0200e120";
		wait for Clk_period;
		Addr <=  "00001100101001";
		Trees_din <= x"05fc1210";
		wait for Clk_period;
		Addr <=  "00001100101010";
		Trees_din <= x"1203ef08";
		wait for Clk_period;
		Addr <=  "00001100101011";
		Trees_din <= x"0f000204";
		wait for Clk_period;
		Addr <=  "00001100101100";
		Trees_din <= x"fffe0d89";
		wait for Clk_period;
		Addr <=  "00001100101101";
		Trees_din <= x"ff660d89";
		wait for Clk_period;
		Addr <=  "00001100101110";
		Trees_din <= x"0e03a004";
		wait for Clk_period;
		Addr <=  "00001100101111";
		Trees_din <= x"ffa20d89";
		wait for Clk_period;
		Addr <=  "00001100110000";
		Trees_din <= x"00c40d89";
		wait for Clk_period;
		Addr <=  "00001100110001";
		Trees_din <= x"04025d08";
		wait for Clk_period;
		Addr <=  "00001100110010";
		Trees_din <= x"0011ff04";
		wait for Clk_period;
		Addr <=  "00001100110011";
		Trees_din <= x"ff7e0d89";
		wait for Clk_period;
		Addr <=  "00001100110100";
		Trees_din <= x"001a0d89";
		wait for Clk_period;
		Addr <=  "00001100110101";
		Trees_din <= x"14013b04";
		wait for Clk_period;
		Addr <=  "00001100110110";
		Trees_din <= x"ffac0d89";
		wait for Clk_period;
		Addr <=  "00001100110111";
		Trees_din <= x"00590d89";
		wait for Clk_period;
		Addr <=  "00001100111000";
		Trees_din <= x"1700210c";
		wait for Clk_period;
		Addr <=  "00001100111001";
		Trees_din <= x"1005bb08";
		wait for Clk_period;
		Addr <=  "00001100111010";
		Trees_din <= x"0a029e04";
		wait for Clk_period;
		Addr <=  "00001100111011";
		Trees_din <= x"ff880d89";
		wait for Clk_period;
		Addr <=  "00001100111100";
		Trees_din <= x"002b0d89";
		wait for Clk_period;
		Addr <=  "00001100111101";
		Trees_din <= x"00eb0d89";
		wait for Clk_period;
		Addr <=  "00001100111110";
		Trees_din <= x"12027b08";
		wait for Clk_period;
		Addr <=  "00001100111111";
		Trees_din <= x"0a01e504";
		wait for Clk_period;
		Addr <=  "00001101000000";
		Trees_din <= x"003c0d89";
		wait for Clk_period;
		Addr <=  "00001101000001";
		Trees_din <= x"ffb00d89";
		wait for Clk_period;
		Addr <=  "00001101000010";
		Trees_din <= x"0e03a004";
		wait for Clk_period;
		Addr <=  "00001101000011";
		Trees_din <= x"00f80d89";
		wait for Clk_period;
		Addr <=  "00001101000100";
		Trees_din <= x"000c0d89";
		wait for Clk_period;
		Addr <=  "00001101000101";
		Trees_din <= x"00192f38";
		wait for Clk_period;
		Addr <=  "00001101000110";
		Trees_din <= x"020e8d20";
		wait for Clk_period;
		Addr <=  "00001101000111";
		Trees_din <= x"08035610";
		wait for Clk_period;
		Addr <=  "00001101001000";
		Trees_din <= x"1e007108";
		wait for Clk_period;
		Addr <=  "00001101001001";
		Trees_din <= x"0e025204";
		wait for Clk_period;
		Addr <=  "00001101001010";
		Trees_din <= x"005b0d89";
		wait for Clk_period;
		Addr <=  "00001101001011";
		Trees_din <= x"00090d89";
		wait for Clk_period;
		Addr <=  "00001101001100";
		Trees_din <= x"03f94d04";
		wait for Clk_period;
		Addr <=  "00001101001101";
		Trees_din <= x"ffd10d89";
		wait for Clk_period;
		Addr <=  "00001101001110";
		Trees_din <= x"002c0d89";
		wait for Clk_period;
		Addr <=  "00001101001111";
		Trees_din <= x"0c02d908";
		wait for Clk_period;
		Addr <=  "00001101010000";
		Trees_din <= x"12fc3904";
		wait for Clk_period;
		Addr <=  "00001101010001";
		Trees_din <= x"008a0d89";
		wait for Clk_period;
		Addr <=  "00001101010010";
		Trees_din <= x"ff770d89";
		wait for Clk_period;
		Addr <=  "00001101010011";
		Trees_din <= x"10028704";
		wait for Clk_period;
		Addr <=  "00001101010100";
		Trees_din <= x"ffc80d89";
		wait for Clk_period;
		Addr <=  "00001101010101";
		Trees_din <= x"00a80d89";
		wait for Clk_period;
		Addr <=  "00001101010110";
		Trees_din <= x"0bf9680c";
		wait for Clk_period;
		Addr <=  "00001101010111";
		Trees_din <= x"0bf95b08";
		wait for Clk_period;
		Addr <=  "00001101011000";
		Trees_din <= x"0f018f04";
		wait for Clk_period;
		Addr <=  "00001101011001";
		Trees_din <= x"00970d89";
		wait for Clk_period;
		Addr <=  "00001101011010";
		Trees_din <= x"ffe20d89";
		wait for Clk_period;
		Addr <=  "00001101011011";
		Trees_din <= x"ff150d89";
		wait for Clk_period;
		Addr <=  "00001101011100";
		Trees_din <= x"010f7408";
		wait for Clk_period;
		Addr <=  "00001101011101";
		Trees_din <= x"00119204";
		wait for Clk_period;
		Addr <=  "00001101011110";
		Trees_din <= x"00980d89";
		wait for Clk_period;
		Addr <=  "00001101011111";
		Trees_din <= x"00070d89";
		wait for Clk_period;
		Addr <=  "00001101100000";
		Trees_din <= x"ffc10d89";
		wait for Clk_period;
		Addr <=  "00001101100001";
		Trees_din <= x"ff710d89";
		wait for Clk_period;
		Addr <=  "00001101100010";
		Trees_din <= x"00167654";
		wait for Clk_period;
		Addr <=  "00001101100011";
		Trees_din <= x"0205be28";
		wait for Clk_period;
		Addr <=  "00001101100100";
		Trees_din <= x"03f84908";
		wait for Clk_period;
		Addr <=  "00001101100101";
		Trees_din <= x"0b056704";
		wait for Clk_period;
		Addr <=  "00001101100110";
		Trees_din <= x"ff6b0e45";
		wait for Clk_period;
		Addr <=  "00001101100111";
		Trees_din <= x"00140e45";
		wait for Clk_period;
		Addr <=  "00001101101000";
		Trees_din <= x"0200e110";
		wait for Clk_period;
		Addr <=  "00001101101001";
		Trees_din <= x"05fc3808";
		wait for Clk_period;
		Addr <=  "00001101101010";
		Trees_din <= x"1203f704";
		wait for Clk_period;
		Addr <=  "00001101101011";
		Trees_din <= x"ff7f0e45";
		wait for Clk_period;
		Addr <=  "00001101101100";
		Trees_din <= x"00280e45";
		wait for Clk_period;
		Addr <=  "00001101101101";
		Trees_din <= x"1e005904";
		wait for Clk_period;
		Addr <=  "00001101101110";
		Trees_din <= x"ff6e0e45";
		wait for Clk_period;
		Addr <=  "00001101101111";
		Trees_din <= x"00140e45";
		wait for Clk_period;
		Addr <=  "00001101110000";
		Trees_din <= x"07005a08";
		wait for Clk_period;
		Addr <=  "00001101110001";
		Trees_din <= x"0d033104";
		wait for Clk_period;
		Addr <=  "00001101110010";
		Trees_din <= x"00350e45";
		wait for Clk_period;
		Addr <=  "00001101110011";
		Trees_din <= x"ffc20e45";
		wait for Clk_period;
		Addr <=  "00001101110100";
		Trees_din <= x"09004804";
		wait for Clk_period;
		Addr <=  "00001101110101";
		Trees_din <= x"00b10e45";
		wait for Clk_period;
		Addr <=  "00001101110110";
		Trees_din <= x"ffa50e45";
		wait for Clk_period;
		Addr <=  "00001101110111";
		Trees_din <= x"0211fd20";
		wait for Clk_period;
		Addr <=  "00001101111000";
		Trees_din <= x"00fde510";
		wait for Clk_period;
		Addr <=  "00001101111001";
		Trees_din <= x"07005508";
		wait for Clk_period;
		Addr <=  "00001101111010";
		Trees_din <= x"04070604";
		wait for Clk_period;
		Addr <=  "00001101111011";
		Trees_din <= x"00910e45";
		wait for Clk_period;
		Addr <=  "00001101111100";
		Trees_din <= x"ff6f0e45";
		wait for Clk_period;
		Addr <=  "00001101111101";
		Trees_din <= x"08028d04";
		wait for Clk_period;
		Addr <=  "00001101111110";
		Trees_din <= x"00d30e45";
		wait for Clk_period;
		Addr <=  "00001101111111";
		Trees_din <= x"00290e45";
		wait for Clk_period;
		Addr <=  "00001110000000";
		Trees_din <= x"10068308";
		wait for Clk_period;
		Addr <=  "00001110000001";
		Trees_din <= x"06f27e04";
		wait for Clk_period;
		Addr <=  "00001110000010";
		Trees_din <= x"ffec0e45";
		wait for Clk_period;
		Addr <=  "00001110000011";
		Trees_din <= x"00300e45";
		wait for Clk_period;
		Addr <=  "00001110000100";
		Trees_din <= x"0f02fb04";
		wait for Clk_period;
		Addr <=  "00001110000101";
		Trees_din <= x"00e30e45";
		wait for Clk_period;
		Addr <=  "00001110000110";
		Trees_din <= x"ffcf0e45";
		wait for Clk_period;
		Addr <=  "00001110000111";
		Trees_din <= x"1d005608";
		wait for Clk_period;
		Addr <=  "00001110001000";
		Trees_din <= x"000fd304";
		wait for Clk_period;
		Addr <=  "00001110001001";
		Trees_din <= x"00a20e45";
		wait for Clk_period;
		Addr <=  "00001110001010";
		Trees_din <= x"fffa0e45";
		wait for Clk_period;
		Addr <=  "00001110001011";
		Trees_din <= x"ffd10e45";
		wait for Clk_period;
		Addr <=  "00001110001100";
		Trees_din <= x"0a07cb08";
		wait for Clk_period;
		Addr <=  "00001110001101";
		Trees_din <= x"0c03f804";
		wait for Clk_period;
		Addr <=  "00001110001110";
		Trees_din <= x"ff670e45";
		wait for Clk_period;
		Addr <=  "00001110001111";
		Trees_din <= x"003a0e45";
		wait for Clk_period;
		Addr <=  "00001110010000";
		Trees_din <= x"00420e45";
		wait for Clk_period;
		Addr <=  "00001110010001";
		Trees_din <= x"0016766c";
		wait for Clk_period;
		Addr <=  "00001110010010";
		Trees_din <= x"0209133c";
		wait for Clk_period;
		Addr <=  "00001110010011";
		Trees_din <= x"02026c20";
		wait for Clk_period;
		Addr <=  "00001110010100";
		Trees_din <= x"10057a10";
		wait for Clk_period;
		Addr <=  "00001110010101";
		Trees_din <= x"21000008";
		wait for Clk_period;
		Addr <=  "00001110010110";
		Trees_din <= x"1203c004";
		wait for Clk_period;
		Addr <=  "00001110010111";
		Trees_din <= x"ffa60f31";
		wait for Clk_period;
		Addr <=  "00001110011000";
		Trees_din <= x"00290f31";
		wait for Clk_period;
		Addr <=  "00001110011001";
		Trees_din <= x"02ffc504";
		wait for Clk_period;
		Addr <=  "00001110011010";
		Trees_din <= x"ff8d0f31";
		wait for Clk_period;
		Addr <=  "00001110011011";
		Trees_din <= x"00ab0f31";
		wait for Clk_period;
		Addr <=  "00001110011100";
		Trees_din <= x"0d024408";
		wait for Clk_period;
		Addr <=  "00001110011101";
		Trees_din <= x"1a008904";
		wait for Clk_period;
		Addr <=  "00001110011110";
		Trees_din <= x"00760f31";
		wait for Clk_period;
		Addr <=  "00001110011111";
		Trees_din <= x"ff790f31";
		wait for Clk_period;
		Addr <=  "00001110100000";
		Trees_din <= x"01074704";
		wait for Clk_period;
		Addr <=  "00001110100001";
		Trees_din <= x"00f70f31";
		wait for Clk_period;
		Addr <=  "00001110100010";
		Trees_din <= x"ffaf0f31";
		wait for Clk_period;
		Addr <=  "00001110100011";
		Trees_din <= x"0f00060c";
		wait for Clk_period;
		Addr <=  "00001110100100";
		Trees_din <= x"17000404";
		wait for Clk_period;
		Addr <=  "00001110100101";
		Trees_din <= x"ff7a0f31";
		wait for Clk_period;
		Addr <=  "00001110100110";
		Trees_din <= x"05f8c104";
		wait for Clk_period;
		Addr <=  "00001110100111";
		Trees_din <= x"ffa30f31";
		wait for Clk_period;
		Addr <=  "00001110101000";
		Trees_din <= x"00a20f31";
		wait for Clk_period;
		Addr <=  "00001110101001";
		Trees_din <= x"14028008";
		wait for Clk_period;
		Addr <=  "00001110101010";
		Trees_din <= x"03f94d04";
		wait for Clk_period;
		Addr <=  "00001110101011";
		Trees_din <= x"ff9c0f31";
		wait for Clk_period;
		Addr <=  "00001110101100";
		Trees_din <= x"fffb0f31";
		wait for Clk_period;
		Addr <=  "00001110101101";
		Trees_din <= x"15009604";
		wait for Clk_period;
		Addr <=  "00001110101110";
		Trees_din <= x"fff20f31";
		wait for Clk_period;
		Addr <=  "00001110101111";
		Trees_din <= x"00720f31";
		wait for Clk_period;
		Addr <=  "00001110110000";
		Trees_din <= x"0c022d18";
		wait for Clk_period;
		Addr <=  "00001110110001";
		Trees_din <= x"1f00000c";
		wait for Clk_period;
		Addr <=  "00001110110010";
		Trees_din <= x"0407e108";
		wait for Clk_period;
		Addr <=  "00001110110011";
		Trees_din <= x"1900a204";
		wait for Clk_period;
		Addr <=  "00001110110100";
		Trees_din <= x"00260f31";
		wait for Clk_period;
		Addr <=  "00001110110101";
		Trees_din <= x"00820f31";
		wait for Clk_period;
		Addr <=  "00001110110110";
		Trees_din <= x"ff700f31";
		wait for Clk_period;
		Addr <=  "00001110110111";
		Trees_din <= x"07004d04";
		wait for Clk_period;
		Addr <=  "00001110111000";
		Trees_din <= x"00770f31";
		wait for Clk_period;
		Addr <=  "00001110111001";
		Trees_din <= x"0d011004";
		wait for Clk_period;
		Addr <=  "00001110111010";
		Trees_din <= x"00210f31";
		wait for Clk_period;
		Addr <=  "00001110111011";
		Trees_din <= x"ff1a0f31";
		wait for Clk_period;
		Addr <=  "00001110111100";
		Trees_din <= x"07005e10";
		wait for Clk_period;
		Addr <=  "00001110111101";
		Trees_din <= x"11048e08";
		wait for Clk_period;
		Addr <=  "00001110111110";
		Trees_din <= x"09005d04";
		wait for Clk_period;
		Addr <=  "00001110111111";
		Trees_din <= x"00800f31";
		wait for Clk_period;
		Addr <=  "00001111000000";
		Trees_din <= x"ffc90f31";
		wait for Clk_period;
		Addr <=  "00001111000001";
		Trees_din <= x"09005404";
		wait for Clk_period;
		Addr <=  "00001111000010";
		Trees_din <= x"005c0f31";
		wait for Clk_period;
		Addr <=  "00001111000011";
		Trees_din <= x"ff6d0f31";
		wait for Clk_period;
		Addr <=  "00001111000100";
		Trees_din <= x"12004604";
		wait for Clk_period;
		Addr <=  "00001111000101";
		Trees_din <= x"00280f31";
		wait for Clk_period;
		Addr <=  "00001111000110";
		Trees_din <= x"ff380f31";
		wait for Clk_period;
		Addr <=  "00001111000111";
		Trees_din <= x"0a07cb08";
		wait for Clk_period;
		Addr <=  "00001111001000";
		Trees_din <= x"0c03f804";
		wait for Clk_period;
		Addr <=  "00001111001001";
		Trees_din <= x"ff680f31";
		wait for Clk_period;
		Addr <=  "00001111001010";
		Trees_din <= x"003a0f31";
		wait for Clk_period;
		Addr <=  "00001111001011";
		Trees_din <= x"003e0f31";
		wait for Clk_period;
		Addr <=  "00001111001100";
		Trees_din <= x"0016764c";
		wait for Clk_period;
		Addr <=  "00001111001101";
		Trees_din <= x"02091320";
		wait for Clk_period;
		Addr <=  "00001111001110";
		Trees_din <= x"02fce404";
		wait for Clk_period;
		Addr <=  "00001111001111";
		Trees_din <= x"ff730fdd";
		wait for Clk_period;
		Addr <=  "00001111010000";
		Trees_din <= x"010f7410";
		wait for Clk_period;
		Addr <=  "00001111010001";
		Trees_din <= x"1104aa08";
		wait for Clk_period;
		Addr <=  "00001111010010";
		Trees_din <= x"08035f04";
		wait for Clk_period;
		Addr <=  "00001111010011";
		Trees_din <= x"000e0fdd";
		wait for Clk_period;
		Addr <=  "00001111010100";
		Trees_din <= x"ffad0fdd";
		wait for Clk_period;
		Addr <=  "00001111010101";
		Trees_din <= x"1b003f04";
		wait for Clk_period;
		Addr <=  "00001111010110";
		Trees_din <= x"ff600fdd";
		wait for Clk_period;
		Addr <=  "00001111010111";
		Trees_din <= x"fff70fdd";
		wait for Clk_period;
		Addr <=  "00001111011000";
		Trees_din <= x"02085c08";
		wait for Clk_period;
		Addr <=  "00001111011001";
		Trees_din <= x"11046804";
		wait for Clk_period;
		Addr <=  "00001111011010";
		Trees_din <= x"ff840fdd";
		wait for Clk_period;
		Addr <=  "00001111011011";
		Trees_din <= x"005a0fdd";
		wait for Clk_period;
		Addr <=  "00001111011100";
		Trees_din <= x"008e0fdd";
		wait for Clk_period;
		Addr <=  "00001111011101";
		Trees_din <= x"0211fd20";
		wait for Clk_period;
		Addr <=  "00001111011110";
		Trees_din <= x"06f2f010";
		wait for Clk_period;
		Addr <=  "00001111011111";
		Trees_din <= x"0c00be08";
		wait for Clk_period;
		Addr <=  "00001111100000";
		Trees_din <= x"09004904";
		wait for Clk_period;
		Addr <=  "00001111100001";
		Trees_din <= x"004d0fdd";
		wait for Clk_period;
		Addr <=  "00001111100010";
		Trees_din <= x"ff680fdd";
		wait for Clk_period;
		Addr <=  "00001111100011";
		Trees_din <= x"0003aa04";
		wait for Clk_period;
		Addr <=  "00001111100100";
		Trees_din <= x"007e0fdd";
		wait for Clk_period;
		Addr <=  "00001111100101";
		Trees_din <= x"ffed0fdd";
		wait for Clk_period;
		Addr <=  "00001111100110";
		Trees_din <= x"0c021208";
		wait for Clk_period;
		Addr <=  "00001111100111";
		Trees_din <= x"0c015d04";
		wait for Clk_period;
		Addr <=  "00001111101000";
		Trees_din <= x"00540fdd";
		wait for Clk_period;
		Addr <=  "00001111101001";
		Trees_din <= x"ffd70fdd";
		wait for Clk_period;
		Addr <=  "00001111101010";
		Trees_din <= x"09004d04";
		wait for Clk_period;
		Addr <=  "00001111101011";
		Trees_din <= x"ff970fdd";
		wait for Clk_period;
		Addr <=  "00001111101100";
		Trees_din <= x"00790fdd";
		wait for Clk_period;
		Addr <=  "00001111101101";
		Trees_din <= x"1d005608";
		wait for Clk_period;
		Addr <=  "00001111101110";
		Trees_din <= x"000fd304";
		wait for Clk_period;
		Addr <=  "00001111101111";
		Trees_din <= x"009c0fdd";
		wait for Clk_period;
		Addr <=  "00001111110000";
		Trees_din <= x"fff50fdd";
		wait for Clk_period;
		Addr <=  "00001111110001";
		Trees_din <= x"ffc70fdd";
		wait for Clk_period;
		Addr <=  "00001111110010";
		Trees_din <= x"0c03f808";
		wait for Clk_period;
		Addr <=  "00001111110011";
		Trees_din <= x"0a07cb04";
		wait for Clk_period;
		Addr <=  "00001111110100";
		Trees_din <= x"ff690fdd";
		wait for Clk_period;
		Addr <=  "00001111110101";
		Trees_din <= x"00380fdd";
		wait for Clk_period;
		Addr <=  "00001111110110";
		Trees_din <= x"003c0fdd";
		wait for Clk_period;
		Addr <=  "00001111110111";
		Trees_din <= x"00192f78";
		wait for Clk_period;
		Addr <=  "00001111111000";
		Trees_din <= x"02026c3c";
		wait for Clk_period;
		Addr <=  "00001111111001";
		Trees_din <= x"10057a20";
		wait for Clk_period;
		Addr <=  "00001111111010";
		Trees_din <= x"09005710";
		wait for Clk_period;
		Addr <=  "00001111111011";
		Trees_din <= x"0402ed08";
		wait for Clk_period;
		Addr <=  "00001111111100";
		Trees_din <= x"19006c04";
		wait for Clk_period;
		Addr <=  "00001111111101";
		Trees_din <= x"008c10d1";
		wait for Clk_period;
		Addr <=  "00001111111110";
		Trees_din <= x"ff6f10d1";
		wait for Clk_period;
		Addr <=  "00001111111111";
		Trees_din <= x"04050404";
		wait for Clk_period;
		Addr <=  "00010000000000";
		Trees_din <= x"006810d1";
		wait for Clk_period;
		Addr <=  "00010000000001";
		Trees_din <= x"ff9f10d1";
		wait for Clk_period;
		Addr <=  "00010000000010";
		Trees_din <= x"1b003408";
		wait for Clk_period;
		Addr <=  "00010000000011";
		Trees_din <= x"18003e04";
		wait for Clk_period;
		Addr <=  "00010000000100";
		Trees_din <= x"ffd210d1";
		wait for Clk_period;
		Addr <=  "00010000000101";
		Trees_din <= x"017d10d1";
		wait for Clk_period;
		Addr <=  "00010000000110";
		Trees_din <= x"00fc3a04";
		wait for Clk_period;
		Addr <=  "00010000000111";
		Trees_din <= x"006710d1";
		wait for Clk_period;
		Addr <=  "00010000001000";
		Trees_din <= x"ffa510d1";
		wait for Clk_period;
		Addr <=  "00010000001001";
		Trees_din <= x"19009210";
		wait for Clk_period;
		Addr <=  "00010000001010";
		Trees_din <= x"0d02b508";
		wait for Clk_period;
		Addr <=  "00010000001011";
		Trees_din <= x"07005704";
		wait for Clk_period;
		Addr <=  "00010000001100";
		Trees_din <= x"006410d1";
		wait for Clk_period;
		Addr <=  "00010000001101";
		Trees_din <= x"ffa810d1";
		wait for Clk_period;
		Addr <=  "00010000001110";
		Trees_din <= x"0c030804";
		wait for Clk_period;
		Addr <=  "00010000001111";
		Trees_din <= x"005a10d1";
		wait for Clk_period;
		Addr <=  "00010000010000";
		Trees_din <= x"015810d1";
		wait for Clk_period;
		Addr <=  "00010000010001";
		Trees_din <= x"1c002a08";
		wait for Clk_period;
		Addr <=  "00010000010010";
		Trees_din <= x"0800ba04";
		wait for Clk_period;
		Addr <=  "00010000010011";
		Trees_din <= x"012610d1";
		wait for Clk_period;
		Addr <=  "00010000010100";
		Trees_din <= x"ffab10d1";
		wait for Clk_period;
		Addr <=  "00010000010101";
		Trees_din <= x"ff7810d1";
		wait for Clk_period;
		Addr <=  "00010000010110";
		Trees_din <= x"020e8d20";
		wait for Clk_period;
		Addr <=  "00010000010111";
		Trees_din <= x"00fd6410";
		wait for Clk_period;
		Addr <=  "00010000011000";
		Trees_din <= x"1500a108";
		wait for Clk_period;
		Addr <=  "00010000011001";
		Trees_din <= x"04f8a504";
		wait for Clk_period;
		Addr <=  "00010000011010";
		Trees_din <= x"ff9d10d1";
		wait for Clk_period;
		Addr <=  "00010000011011";
		Trees_din <= x"009e10d1";
		wait for Clk_period;
		Addr <=  "00010000011100";
		Trees_din <= x"04070604";
		wait for Clk_period;
		Addr <=  "00010000011101";
		Trees_din <= x"003c10d1";
		wait for Clk_period;
		Addr <=  "00010000011110";
		Trees_din <= x"ff7310d1";
		wait for Clk_period;
		Addr <=  "00010000011111";
		Trees_din <= x"18004208";
		wait for Clk_period;
		Addr <=  "00010000100000";
		Trees_din <= x"14028004";
		wait for Clk_period;
		Addr <=  "00010000100001";
		Trees_din <= x"000b10d1";
		wait for Clk_period;
		Addr <=  "00010000100010";
		Trees_din <= x"006610d1";
		wait for Clk_period;
		Addr <=  "00010000100011";
		Trees_din <= x"15008f04";
		wait for Clk_period;
		Addr <=  "00010000100100";
		Trees_din <= x"001010d1";
		wait for Clk_period;
		Addr <=  "00010000100101";
		Trees_din <= x"ffcb10d1";
		wait for Clk_period;
		Addr <=  "00010000100110";
		Trees_din <= x"0afb310c";
		wait for Clk_period;
		Addr <=  "00010000100111";
		Trees_din <= x"1102f108";
		wait for Clk_period;
		Addr <=  "00010000101000";
		Trees_din <= x"11007904";
		wait for Clk_period;
		Addr <=  "00010000101001";
		Trees_din <= x"ff6e10d1";
		wait for Clk_period;
		Addr <=  "00010000101010";
		Trees_din <= x"006310d1";
		wait for Clk_period;
		Addr <=  "00010000101011";
		Trees_din <= x"ff4410d1";
		wait for Clk_period;
		Addr <=  "00010000101100";
		Trees_din <= x"1b002c08";
		wait for Clk_period;
		Addr <=  "00010000101101";
		Trees_din <= x"1f000004";
		wait for Clk_period;
		Addr <=  "00010000101110";
		Trees_din <= x"004c10d1";
		wait for Clk_period;
		Addr <=  "00010000101111";
		Trees_din <= x"ff6d10d1";
		wait for Clk_period;
		Addr <=  "00010000110000";
		Trees_din <= x"000fd304";
		wait for Clk_period;
		Addr <=  "00010000110001";
		Trees_din <= x"009d10d1";
		wait for Clk_period;
		Addr <=  "00010000110010";
		Trees_din <= x"001610d1";
		wait for Clk_period;
		Addr <=  "00010000110011";
		Trees_din <= x"ff6b10d1";
		wait for Clk_period;
		Addr <=  "00010000110100";
		Trees_din <= x"00192f64";
		wait for Clk_period;
		Addr <=  "00010000110101";
		Trees_din <= x"02047538";
		wait for Clk_period;
		Addr <=  "00010000110110";
		Trees_din <= x"04022418";
		wait for Clk_period;
		Addr <=  "00010000110111";
		Trees_din <= x"21000110";
		wait for Clk_period;
		Addr <=  "00010000111000";
		Trees_din <= x"08021408";
		wait for Clk_period;
		Addr <=  "00010000111001";
		Trees_din <= x"03fc7704";
		wait for Clk_period;
		Addr <=  "00010000111010";
		Trees_din <= x"ff74119d";
		wait for Clk_period;
		Addr <=  "00010000111011";
		Trees_din <= x"ffcd119d";
		wait for Clk_period;
		Addr <=  "00010000111100";
		Trees_din <= x"0d00cc04";
		wait for Clk_period;
		Addr <=  "00010000111101";
		Trees_din <= x"ff76119d";
		wait for Clk_period;
		Addr <=  "00010000111110";
		Trees_din <= x"0051119d";
		wait for Clk_period;
		Addr <=  "00010000111111";
		Trees_din <= x"07005504";
		wait for Clk_period;
		Addr <=  "00010001000000";
		Trees_din <= x"00de119d";
		wait for Clk_period;
		Addr <=  "00010001000001";
		Trees_din <= x"fffa119d";
		wait for Clk_period;
		Addr <=  "00010001000010";
		Trees_din <= x"0406be10";
		wait for Clk_period;
		Addr <=  "00010001000011";
		Trees_din <= x"0e01da08";
		wait for Clk_period;
		Addr <=  "00010001000100";
		Trees_din <= x"05fc3804";
		wait for Clk_period;
		Addr <=  "00010001000101";
		Trees_din <= x"0012119d";
		wait for Clk_period;
		Addr <=  "00010001000110";
		Trees_din <= x"00a4119d";
		wait for Clk_period;
		Addr <=  "00010001000111";
		Trees_din <= x"01099e04";
		wait for Clk_period;
		Addr <=  "00010001001000";
		Trees_din <= x"ffa9119d";
		wait for Clk_period;
		Addr <=  "00010001001001";
		Trees_din <= x"0088119d";
		wait for Clk_period;
		Addr <=  "00010001001010";
		Trees_din <= x"1101f308";
		wait for Clk_period;
		Addr <=  "00010001001011";
		Trees_din <= x"12fd6804";
		wait for Clk_period;
		Addr <=  "00010001001100";
		Trees_din <= x"0022119d";
		wait for Clk_period;
		Addr <=  "00010001001101";
		Trees_din <= x"ff6f119d";
		wait for Clk_period;
		Addr <=  "00010001001110";
		Trees_din <= x"07005704";
		wait for Clk_period;
		Addr <=  "00010001001111";
		Trees_din <= x"ffa6119d";
		wait for Clk_period;
		Addr <=  "00010001010000";
		Trees_din <= x"004e119d";
		wait for Clk_period;
		Addr <=  "00010001010001";
		Trees_din <= x"0211fd20";
		wait for Clk_period;
		Addr <=  "00010001010010";
		Trees_din <= x"08034310";
		wait for Clk_period;
		Addr <=  "00010001010011";
		Trees_din <= x"0e041108";
		wait for Clk_period;
		Addr <=  "00010001010100";
		Trees_din <= x"0800b204";
		wait for Clk_period;
		Addr <=  "00010001010101";
		Trees_din <= x"0009119d";
		wait for Clk_period;
		Addr <=  "00010001010110";
		Trees_din <= x"0038119d";
		wait for Clk_period;
		Addr <=  "00010001010111";
		Trees_din <= x"10fade04";
		wait for Clk_period;
		Addr <=  "00010001011000";
		Trees_din <= x"005a119d";
		wait for Clk_period;
		Addr <=  "00010001011001";
		Trees_din <= x"ff86119d";
		wait for Clk_period;
		Addr <=  "00010001011010";
		Trees_din <= x"0d011008";
		wait for Clk_period;
		Addr <=  "00010001011011";
		Trees_din <= x"17000004";
		wait for Clk_period;
		Addr <=  "00010001011100";
		Trees_din <= x"ff78119d";
		wait for Clk_period;
		Addr <=  "00010001011101";
		Trees_din <= x"0042119d";
		wait for Clk_period;
		Addr <=  "00010001011110";
		Trees_din <= x"18003b04";
		wait for Clk_period;
		Addr <=  "00010001011111";
		Trees_din <= x"ff23119d";
		wait for Clk_period;
		Addr <=  "00010001100000";
		Trees_din <= x"ffd4119d";
		wait for Clk_period;
		Addr <=  "00010001100001";
		Trees_din <= x"1a008e04";
		wait for Clk_period;
		Addr <=  "00010001100010";
		Trees_din <= x"ffbc119d";
		wait for Clk_period;
		Addr <=  "00010001100011";
		Trees_din <= x"000fd304";
		wait for Clk_period;
		Addr <=  "00010001100100";
		Trees_din <= x"0097119d";
		wait for Clk_period;
		Addr <=  "00010001100101";
		Trees_din <= x"fff4119d";
		wait for Clk_period;
		Addr <=  "00010001100110";
		Trees_din <= x"ff6d119d";
		wait for Clk_period;
		Addr <=  "00010001100111";
		Trees_din <= x"00192f60";
		wait for Clk_period;
		Addr <=  "00010001101000";
		Trees_din <= x"02026c34";
		wait for Clk_period;
		Addr <=  "00010001101001";
		Trees_din <= x"1005661c";
		wait for Clk_period;
		Addr <=  "00010001101010";
		Trees_din <= x"0900570c";
		wait for Clk_period;
		Addr <=  "00010001101011";
		Trees_din <= x"19007104";
		wait for Clk_period;
		Addr <=  "00010001101100";
		Trees_din <= x"007e1261";
		wait for Clk_period;
		Addr <=  "00010001101101";
		Trees_din <= x"0402ed04";
		wait for Clk_period;
		Addr <=  "00010001101110";
		Trees_din <= x"ff751261";
		wait for Clk_period;
		Addr <=  "00010001101111";
		Trees_din <= x"ffda1261";
		wait for Clk_period;
		Addr <=  "00010001110000";
		Trees_din <= x"07005908";
		wait for Clk_period;
		Addr <=  "00010001110001";
		Trees_din <= x"02fece04";
		wait for Clk_period;
		Addr <=  "00010001110010";
		Trees_din <= x"ff861261";
		wait for Clk_period;
		Addr <=  "00010001110011";
		Trees_din <= x"006a1261";
		wait for Clk_period;
		Addr <=  "00010001110100";
		Trees_din <= x"00f9b904";
		wait for Clk_period;
		Addr <=  "00010001110101";
		Trees_din <= x"004e1261";
		wait for Clk_period;
		Addr <=  "00010001110110";
		Trees_din <= x"ff871261";
		wait for Clk_period;
		Addr <=  "00010001110111";
		Trees_din <= x"1900920c";
		wait for Clk_period;
		Addr <=  "00010001111000";
		Trees_din <= x"0d013f04";
		wait for Clk_period;
		Addr <=  "00010001111001";
		Trees_din <= x"fff21261";
		wait for Clk_period;
		Addr <=  "00010001111010";
		Trees_din <= x"17000004";
		wait for Clk_period;
		Addr <=  "00010001111011";
		Trees_din <= x"01071261";
		wait for Clk_period;
		Addr <=  "00010001111100";
		Trees_din <= x"00261261";
		wait for Clk_period;
		Addr <=  "00010001111101";
		Trees_din <= x"0800ba08";
		wait for Clk_period;
		Addr <=  "00010001111110";
		Trees_din <= x"1900a604";
		wait for Clk_period;
		Addr <=  "00010001111111";
		Trees_din <= x"ffaf1261";
		wait for Clk_period;
		Addr <=  "00010010000000";
		Trees_din <= x"00f41261";
		wait for Clk_period;
		Addr <=  "00010010000001";
		Trees_din <= x"ff7b1261";
		wait for Clk_period;
		Addr <=  "00010010000010";
		Trees_din <= x"0211fd20";
		wait for Clk_period;
		Addr <=  "00010010000011";
		Trees_din <= x"00fd6410";
		wait for Clk_period;
		Addr <=  "00010010000100";
		Trees_din <= x"1500a108";
		wait for Clk_period;
		Addr <=  "00010010000101";
		Trees_din <= x"05fc1d04";
		wait for Clk_period;
		Addr <=  "00010010000110";
		Trees_din <= x"00a31261";
		wait for Clk_period;
		Addr <=  "00010010000111";
		Trees_din <= x"fff71261";
		wait for Clk_period;
		Addr <=  "00010010001000";
		Trees_din <= x"01fe1204";
		wait for Clk_period;
		Addr <=  "00010010001001";
		Trees_din <= x"00891261";
		wait for Clk_period;
		Addr <=  "00010010001010";
		Trees_din <= x"ffb71261";
		wait for Clk_period;
		Addr <=  "00010010001011";
		Trees_din <= x"1d004308";
		wait for Clk_period;
		Addr <=  "00010010001100";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00010010001101";
		Trees_din <= x"000c1261";
		wait for Clk_period;
		Addr <=  "00010010001110";
		Trees_din <= x"00811261";
		wait for Clk_period;
		Addr <=  "00010010001111";
		Trees_din <= x"07005e04";
		wait for Clk_period;
		Addr <=  "00010010010000";
		Trees_din <= x"00011261";
		wait for Clk_period;
		Addr <=  "00010010010001";
		Trees_din <= x"ff5f1261";
		wait for Clk_period;
		Addr <=  "00010010010010";
		Trees_din <= x"1a008e04";
		wait for Clk_period;
		Addr <=  "00010010010011";
		Trees_din <= x"ffbe1261";
		wait for Clk_period;
		Addr <=  "00010010010100";
		Trees_din <= x"000fd304";
		wait for Clk_period;
		Addr <=  "00010010010101";
		Trees_din <= x"00931261";
		wait for Clk_period;
		Addr <=  "00010010010110";
		Trees_din <= x"fff81261";
		wait for Clk_period;
		Addr <=  "00010010010111";
		Trees_din <= x"ff6f1261";
		wait for Clk_period;
		Addr <=  "00010010011000";
		Trees_din <= x"00192f30";
		wait for Clk_period;
		Addr <=  "00010010011001";
		Trees_din <= x"02fce404";
		wait for Clk_period;
		Addr <=  "00010010011010";
		Trees_din <= x"ff7a12c5";
		wait for Clk_period;
		Addr <=  "00010010011011";
		Trees_din <= x"0211fd20";
		wait for Clk_period;
		Addr <=  "00010010011100";
		Trees_din <= x"00fc3a10";
		wait for Clk_period;
		Addr <=  "00010010011101";
		Trees_din <= x"0405b608";
		wait for Clk_period;
		Addr <=  "00010010011110";
		Trees_din <= x"04fe8104";
		wait for Clk_period;
		Addr <=  "00010010011111";
		Trees_din <= x"ffe512c5";
		wait for Clk_period;
		Addr <=  "00010010100000";
		Trees_din <= x"00ae12c5";
		wait for Clk_period;
		Addr <=  "00010010100001";
		Trees_din <= x"1203c004";
		wait for Clk_period;
		Addr <=  "00010010100010";
		Trees_din <= x"ffde12c5";
		wait for Clk_period;
		Addr <=  "00010010100011";
		Trees_din <= x"007d12c5";
		wait for Clk_period;
		Addr <=  "00010010100100";
		Trees_din <= x"02047508";
		wait for Clk_period;
		Addr <=  "00010010100101";
		Trees_din <= x"1500a604";
		wait for Clk_period;
		Addr <=  "00010010100110";
		Trees_din <= x"ffd912c5";
		wait for Clk_period;
		Addr <=  "00010010100111";
		Trees_din <= x"002912c5";
		wait for Clk_period;
		Addr <=  "00010010101000";
		Trees_din <= x"0e025a04";
		wait for Clk_period;
		Addr <=  "00010010101001";
		Trees_din <= x"001b12c5";
		wait for Clk_period;
		Addr <=  "00010010101010";
		Trees_din <= x"ffec12c5";
		wait for Clk_period;
		Addr <=  "00010010101011";
		Trees_din <= x"1a008e04";
		wait for Clk_period;
		Addr <=  "00010010101100";
		Trees_din <= x"ffc312c5";
		wait for Clk_period;
		Addr <=  "00010010101101";
		Trees_din <= x"000fd304";
		wait for Clk_period;
		Addr <=  "00010010101110";
		Trees_din <= x"009012c5";
		wait for Clk_period;
		Addr <=  "00010010101111";
		Trees_din <= x"fff912c5";
		wait for Clk_period;
		Addr <=  "00010010110000";
		Trees_din <= x"ff7212c5";
		wait for Clk_period;
		Addr <=  "00010010110001";
		Trees_din <= x"00192f30";
		wait for Clk_period;
		Addr <=  "00010010110010";
		Trees_din <= x"02fce404";
		wait for Clk_period;
		Addr <=  "00010010110011";
		Trees_din <= x"ff7e1329";
		wait for Clk_period;
		Addr <=  "00010010110100";
		Trees_din <= x"0211fd20";
		wait for Clk_period;
		Addr <=  "00010010110101";
		Trees_din <= x"08036910";
		wait for Clk_period;
		Addr <=  "00010010110110";
		Trees_din <= x"1104aa08";
		wait for Clk_period;
		Addr <=  "00010010110111";
		Trees_din <= x"08020d04";
		wait for Clk_period;
		Addr <=  "00010010111000";
		Trees_din <= x"00061329";
		wait for Clk_period;
		Addr <=  "00010010111001";
		Trees_din <= x"002e1329";
		wait for Clk_period;
		Addr <=  "00010010111010";
		Trees_din <= x"020cbe04";
		wait for Clk_period;
		Addr <=  "00010010111011";
		Trees_din <= x"ff821329";
		wait for Clk_period;
		Addr <=  "00010010111100";
		Trees_din <= x"00441329";
		wait for Clk_period;
		Addr <=  "00010010111101";
		Trees_din <= x"0c02ba08";
		wait for Clk_period;
		Addr <=  "00010010111110";
		Trees_din <= x"09004d04";
		wait for Clk_period;
		Addr <=  "00010010111111";
		Trees_din <= x"005b1329";
		wait for Clk_period;
		Addr <=  "00010011000000";
		Trees_din <= x"ff721329";
		wait for Clk_period;
		Addr <=  "00010011000001";
		Trees_din <= x"11028704";
		wait for Clk_period;
		Addr <=  "00010011000010";
		Trees_din <= x"ffc11329";
		wait for Clk_period;
		Addr <=  "00010011000011";
		Trees_din <= x"00e01329";
		wait for Clk_period;
		Addr <=  "00010011000100";
		Trees_din <= x"1a008e04";
		wait for Clk_period;
		Addr <=  "00010011000101";
		Trees_din <= x"ffc71329";
		wait for Clk_period;
		Addr <=  "00010011000110";
		Trees_din <= x"000fd304";
		wait for Clk_period;
		Addr <=  "00010011000111";
		Trees_din <= x"008d1329";
		wait for Clk_period;
		Addr <=  "00010011001000";
		Trees_din <= x"fff71329";
		wait for Clk_period;
		Addr <=  "00010011001001";
		Trees_din <= x"ff751329";
		wait for Clk_period;
		Addr <=  "00010011001010";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00010011001011";
		Trees_din <= x"00192f64";
		wait for Clk_period;
		Addr <=  "00010011001100";
		Trees_din <= x"0209132c";
		wait for Clk_period;
		Addr <=  "00010011001101";
		Trees_din <= x"13f86f0c";
		wait for Clk_period;
		Addr <=  "00010011001110";
		Trees_din <= x"1403bd08";
		wait for Clk_period;
		Addr <=  "00010011001111";
		Trees_din <= x"1900a204";
		wait for Clk_period;
		Addr <=  "00010011010000";
		Trees_din <= x"ff6113f9";
		wait for Clk_period;
		Addr <=  "00010011010001";
		Trees_din <= x"ffdc13f9";
		wait for Clk_period;
		Addr <=  "00010011010010";
		Trees_din <= x"008713f9";
		wait for Clk_period;
		Addr <=  "00010011010011";
		Trees_din <= x"1702f910";
		wait for Clk_period;
		Addr <=  "00010011010100";
		Trees_din <= x"1400c308";
		wait for Clk_period;
		Addr <=  "00010011010101";
		Trees_din <= x"04ff5704";
		wait for Clk_period;
		Addr <=  "00010011010110";
		Trees_din <= x"fffb13f9";
		wait for Clk_period;
		Addr <=  "00010011010111";
		Trees_din <= x"ff8113f9";
		wait for Clk_period;
		Addr <=  "00010011011000";
		Trees_din <= x"1a00e004";
		wait for Clk_period;
		Addr <=  "00010011011001";
		Trees_din <= x"001113f9";
		wait for Clk_period;
		Addr <=  "00010011011010";
		Trees_din <= x"ffda13f9";
		wait for Clk_period;
		Addr <=  "00010011011011";
		Trees_din <= x"0f000608";
		wait for Clk_period;
		Addr <=  "00010011011100";
		Trees_din <= x"19009904";
		wait for Clk_period;
		Addr <=  "00010011011101";
		Trees_din <= x"002313f9";
		wait for Clk_period;
		Addr <=  "00010011011110";
		Trees_din <= x"010c13f9";
		wait for Clk_period;
		Addr <=  "00010011011111";
		Trees_din <= x"04004504";
		wait for Clk_period;
		Addr <=  "00010011100000";
		Trees_din <= x"ffb313f9";
		wait for Clk_period;
		Addr <=  "00010011100001";
		Trees_din <= x"004c13f9";
		wait for Clk_period;
		Addr <=  "00010011100010";
		Trees_din <= x"0c022d20";
		wait for Clk_period;
		Addr <=  "00010011100011";
		Trees_din <= x"08028d10";
		wait for Clk_period;
		Addr <=  "00010011100100";
		Trees_din <= x"0801cf08";
		wait for Clk_period;
		Addr <=  "00010011100101";
		Trees_din <= x"06f19b04";
		wait for Clk_period;
		Addr <=  "00010011100110";
		Trees_din <= x"ffb813f9";
		wait for Clk_period;
		Addr <=  "00010011100111";
		Trees_din <= x"001813f9";
		wait for Clk_period;
		Addr <=  "00010011101000";
		Trees_din <= x"08024c04";
		wait for Clk_period;
		Addr <=  "00010011101001";
		Trees_din <= x"00ab13f9";
		wait for Clk_period;
		Addr <=  "00010011101010";
		Trees_din <= x"001d13f9";
		wait for Clk_period;
		Addr <=  "00010011101011";
		Trees_din <= x"0d00dd08";
		wait for Clk_period;
		Addr <=  "00010011101100";
		Trees_din <= x"0f017304";
		wait for Clk_period;
		Addr <=  "00010011101101";
		Trees_din <= x"008213f9";
		wait for Clk_period;
		Addr <=  "00010011101110";
		Trees_din <= x"ff9f13f9";
		wait for Clk_period;
		Addr <=  "00010011101111";
		Trees_din <= x"13ff4404";
		wait for Clk_period;
		Addr <=  "00010011110000";
		Trees_din <= x"ffd213f9";
		wait for Clk_period;
		Addr <=  "00010011110001";
		Trees_din <= x"ff1413f9";
		wait for Clk_period;
		Addr <=  "00010011110010";
		Trees_din <= x"07005e10";
		wait for Clk_period;
		Addr <=  "00010011110011";
		Trees_din <= x"09004c08";
		wait for Clk_period;
		Addr <=  "00010011110100";
		Trees_din <= x"00050804";
		wait for Clk_period;
		Addr <=  "00010011110101";
		Trees_din <= x"005513f9";
		wait for Clk_period;
		Addr <=  "00010011110110";
		Trees_din <= x"ff6513f9";
		wait for Clk_period;
		Addr <=  "00010011110111";
		Trees_din <= x"12027d04";
		wait for Clk_period;
		Addr <=  "00010011111000";
		Trees_din <= x"007013f9";
		wait for Clk_period;
		Addr <=  "00010011111001";
		Trees_din <= x"001313f9";
		wait for Clk_period;
		Addr <=  "00010011111010";
		Trees_din <= x"12004604";
		wait for Clk_period;
		Addr <=  "00010011111011";
		Trees_din <= x"000c13f9";
		wait for Clk_period;
		Addr <=  "00010011111100";
		Trees_din <= x"ff4e13f9";
		wait for Clk_period;
		Addr <=  "00010011111101";
		Trees_din <= x"ff7913f9";
		wait for Clk_period;
		Addr <=  "00010011111110";
		Trees_din <= x"00192f38";
		wait for Clk_period;
		Addr <=  "00010011111111";
		Trees_din <= x"02fce404";
		wait for Clk_period;
		Addr <=  "00010100000000";
		Trees_din <= x"ff83146d";
		wait for Clk_period;
		Addr <=  "00010100000001";
		Trees_din <= x"020baf20";
		wait for Clk_period;
		Addr <=  "00010100000010";
		Trees_din <= x"04f95810";
		wait for Clk_period;
		Addr <=  "00010100000011";
		Trees_din <= x"10f97c08";
		wait for Clk_period;
		Addr <=  "00010100000100";
		Trees_din <= x"1a00df04";
		wait for Clk_period;
		Addr <=  "00010100000101";
		Trees_din <= x"ff5c146d";
		wait for Clk_period;
		Addr <=  "00010100000110";
		Trees_din <= x"ffd4146d";
		wait for Clk_period;
		Addr <=  "00010100000111";
		Trees_din <= x"06f64e04";
		wait for Clk_period;
		Addr <=  "00010100001000";
		Trees_din <= x"ffa5146d";
		wait for Clk_period;
		Addr <=  "00010100001001";
		Trees_din <= x"0007146d";
		wait for Clk_period;
		Addr <=  "00010100001010";
		Trees_din <= x"04f9a008";
		wait for Clk_period;
		Addr <=  "00010100001011";
		Trees_din <= x"0e008204";
		wait for Clk_period;
		Addr <=  "00010100001100";
		Trees_din <= x"fff3146d";
		wait for Clk_period;
		Addr <=  "00010100001101";
		Trees_din <= x"00bc146d";
		wait for Clk_period;
		Addr <=  "00010100001110";
		Trees_din <= x"08001504";
		wait for Clk_period;
		Addr <=  "00010100001111";
		Trees_din <= x"ffd4146d";
		wait for Clk_period;
		Addr <=  "00010100010000";
		Trees_din <= x"000d146d";
		wait for Clk_period;
		Addr <=  "00010100010001";
		Trees_din <= x"0001c404";
		wait for Clk_period;
		Addr <=  "00010100010010";
		Trees_din <= x"0091146d";
		wait for Clk_period;
		Addr <=  "00010100010011";
		Trees_din <= x"12012808";
		wait for Clk_period;
		Addr <=  "00010100010100";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00010100010101";
		Trees_din <= x"ffc8146d";
		wait for Clk_period;
		Addr <=  "00010100010110";
		Trees_din <= x"005f146d";
		wait for Clk_period;
		Addr <=  "00010100010111";
		Trees_din <= x"13ff9a04";
		wait for Clk_period;
		Addr <=  "00010100011000";
		Trees_din <= x"ff9d146d";
		wait for Clk_period;
		Addr <=  "00010100011001";
		Trees_din <= x"002d146d";
		wait for Clk_period;
		Addr <=  "00010100011010";
		Trees_din <= x"ff7d146d";
		wait for Clk_period;
		Addr <=  "00010100011011";
		Trees_din <= x"00192f68";
		wait for Clk_period;
		Addr <=  "00010100011100";
		Trees_din <= x"0406be3c";
		wait for Clk_period;
		Addr <=  "00010100011101";
		Trees_din <= x"00fce81c";
		wait for Clk_period;
		Addr <=  "00010100011110";
		Trees_din <= x"1201fc0c";
		wait for Clk_period;
		Addr <=  "00010100011111";
		Trees_din <= x"04fe8104";
		wait for Clk_period;
		Addr <=  "00010100100000";
		Trees_din <= x"ffe01541";
		wait for Clk_period;
		Addr <=  "00010100100001";
		Trees_din <= x"030a7404";
		wait for Clk_period;
		Addr <=  "00010100100010";
		Trees_din <= x"00c51541";
		wait for Clk_period;
		Addr <=  "00010100100011";
		Trees_din <= x"fff21541";
		wait for Clk_period;
		Addr <=  "00010100100100";
		Trees_din <= x"1c003c08";
		wait for Clk_period;
		Addr <=  "00010100100101";
		Trees_din <= x"1500a604";
		wait for Clk_period;
		Addr <=  "00010100100110";
		Trees_din <= x"ff911541";
		wait for Clk_period;
		Addr <=  "00010100100111";
		Trees_din <= x"ffe91541";
		wait for Clk_period;
		Addr <=  "00010100101000";
		Trees_din <= x"01fc0b04";
		wait for Clk_period;
		Addr <=  "00010100101001";
		Trees_din <= x"00821541";
		wait for Clk_period;
		Addr <=  "00010100101010";
		Trees_din <= x"00101541";
		wait for Clk_period;
		Addr <=  "00010100101011";
		Trees_din <= x"1500aa10";
		wait for Clk_period;
		Addr <=  "00010100101100";
		Trees_din <= x"1400dd08";
		wait for Clk_period;
		Addr <=  "00010100101101";
		Trees_din <= x"0b04d704";
		wait for Clk_period;
		Addr <=  "00010100101110";
		Trees_din <= x"ffcd1541";
		wait for Clk_period;
		Addr <=  "00010100101111";
		Trees_din <= x"00311541";
		wait for Clk_period;
		Addr <=  "00010100110000";
		Trees_din <= x"09004d04";
		wait for Clk_period;
		Addr <=  "00010100110001";
		Trees_din <= x"ff9e1541";
		wait for Clk_period;
		Addr <=  "00010100110010";
		Trees_din <= x"00141541";
		wait for Clk_period;
		Addr <=  "00010100110011";
		Trees_din <= x"1d003d08";
		wait for Clk_period;
		Addr <=  "00010100110100";
		Trees_din <= x"08009b04";
		wait for Clk_period;
		Addr <=  "00010100110101";
		Trees_din <= x"00701541";
		wait for Clk_period;
		Addr <=  "00010100110110";
		Trees_din <= x"ffcd1541";
		wait for Clk_period;
		Addr <=  "00010100110111";
		Trees_din <= x"04fb0604";
		wait for Clk_period;
		Addr <=  "00010100111000";
		Trees_din <= x"00421541";
		wait for Clk_period;
		Addr <=  "00010100111001";
		Trees_din <= x"01371541";
		wait for Clk_period;
		Addr <=  "00010100111010";
		Trees_din <= x"09005818";
		wait for Clk_period;
		Addr <=  "00010100111011";
		Trees_din <= x"1b004e10";
		wait for Clk_period;
		Addr <=  "00010100111100";
		Trees_din <= x"06f40308";
		wait for Clk_period;
		Addr <=  "00010100111101";
		Trees_din <= x"1c002e04";
		wait for Clk_period;
		Addr <=  "00010100111110";
		Trees_din <= x"ff541541";
		wait for Clk_period;
		Addr <=  "00010100111111";
		Trees_din <= x"00251541";
		wait for Clk_period;
		Addr <=  "00010101000000";
		Trees_din <= x"1500ac04";
		wait for Clk_period;
		Addr <=  "00010101000001";
		Trees_din <= x"ff5c1541";
		wait for Clk_period;
		Addr <=  "00010101000010";
		Trees_din <= x"ffeb1541";
		wait for Clk_period;
		Addr <=  "00010101000011";
		Trees_din <= x"03008e04";
		wait for Clk_period;
		Addr <=  "00010101000100";
		Trees_din <= x"009a1541";
		wait for Clk_period;
		Addr <=  "00010101000101";
		Trees_din <= x"fff11541";
		wait for Clk_period;
		Addr <=  "00010101000110";
		Trees_din <= x"1d004508";
		wait for Clk_period;
		Addr <=  "00010101000111";
		Trees_din <= x"19009e04";
		wait for Clk_period;
		Addr <=  "00010101001000";
		Trees_din <= x"ff701541";
		wait for Clk_period;
		Addr <=  "00010101001001";
		Trees_din <= x"ffe51541";
		wait for Clk_period;
		Addr <=  "00010101001010";
		Trees_din <= x"1100c904";
		wait for Clk_period;
		Addr <=  "00010101001011";
		Trees_din <= x"ffd21541";
		wait for Clk_period;
		Addr <=  "00010101001100";
		Trees_din <= x"15008b04";
		wait for Clk_period;
		Addr <=  "00010101001101";
		Trees_din <= x"00381541";
		wait for Clk_period;
		Addr <=  "00010101001110";
		Trees_din <= x"00d51541";
		wait for Clk_period;
		Addr <=  "00010101001111";
		Trees_din <= x"ff831541";
		wait for Clk_period;
		Addr <=  "00010101010000";
		Trees_din <= x"0200e140";
		wait for Clk_period;
		Addr <=  "00010101010001";
		Trees_din <= x"05fc1210";
		wait for Clk_period;
		Addr <=  "00010101010010";
		Trees_din <= x"0d027a04";
		wait for Clk_period;
		Addr <=  "00010101010011";
		Trees_din <= x"ff6f1635";
		wait for Clk_period;
		Addr <=  "00010101010100";
		Trees_din <= x"0801f408";
		wait for Clk_period;
		Addr <=  "00010101010101";
		Trees_din <= x"15008204";
		wait for Clk_period;
		Addr <=  "00010101010110";
		Trees_din <= x"006b1635";
		wait for Clk_period;
		Addr <=  "00010101010111";
		Trees_din <= x"ff7d1635";
		wait for Clk_period;
		Addr <=  "00010101011000";
		Trees_din <= x"00c41635";
		wait for Clk_period;
		Addr <=  "00010101011001";
		Trees_din <= x"17002f18";
		wait for Clk_period;
		Addr <=  "00010101011010";
		Trees_din <= x"07005708";
		wait for Clk_period;
		Addr <=  "00010101011011";
		Trees_din <= x"12fda004";
		wait for Clk_period;
		Addr <=  "00010101011100";
		Trees_din <= x"001c1635";
		wait for Clk_period;
		Addr <=  "00010101011101";
		Trees_din <= x"ff841635";
		wait for Clk_period;
		Addr <=  "00010101011110";
		Trees_din <= x"13ff5808";
		wait for Clk_period;
		Addr <=  "00010101011111";
		Trees_din <= x"1402b804";
		wait for Clk_period;
		Addr <=  "00010101100000";
		Trees_din <= x"01221635";
		wait for Clk_period;
		Addr <=  "00010101100001";
		Trees_din <= x"001e1635";
		wait for Clk_period;
		Addr <=  "00010101100010";
		Trees_din <= x"06f57204";
		wait for Clk_period;
		Addr <=  "00010101100011";
		Trees_din <= x"00901635";
		wait for Clk_period;
		Addr <=  "00010101100100";
		Trees_din <= x"ff881635";
		wait for Clk_period;
		Addr <=  "00010101100101";
		Trees_din <= x"0b04dc10";
		wait for Clk_period;
		Addr <=  "00010101100110";
		Trees_din <= x"0bf95b08";
		wait for Clk_period;
		Addr <=  "00010101100111";
		Trees_din <= x"00005104";
		wait for Clk_period;
		Addr <=  "00010101101000";
		Trees_din <= x"00b01635";
		wait for Clk_period;
		Addr <=  "00010101101001";
		Trees_din <= x"ffa71635";
		wait for Clk_period;
		Addr <=  "00010101101010";
		Trees_din <= x"0f029904";
		wait for Clk_period;
		Addr <=  "00010101101011";
		Trees_din <= x"ff6c1635";
		wait for Clk_period;
		Addr <=  "00010101101100";
		Trees_din <= x"fffc1635";
		wait for Clk_period;
		Addr <=  "00010101101101";
		Trees_din <= x"0d019e04";
		wait for Clk_period;
		Addr <=  "00010101101110";
		Trees_din <= x"00a21635";
		wait for Clk_period;
		Addr <=  "00010101101111";
		Trees_din <= x"00061635";
		wait for Clk_period;
		Addr <=  "00010101110000";
		Trees_din <= x"21000128";
		wait for Clk_period;
		Addr <=  "00010101110001";
		Trees_din <= x"01fb5b10";
		wait for Clk_period;
		Addr <=  "00010101110010";
		Trees_din <= x"0e01e30c";
		wait for Clk_period;
		Addr <=  "00010101110011";
		Trees_din <= x"16017504";
		wait for Clk_period;
		Addr <=  "00010101110100";
		Trees_din <= x"00de1635";
		wait for Clk_period;
		Addr <=  "00010101110101";
		Trees_din <= x"0c00ed04";
		wait for Clk_period;
		Addr <=  "00010101110110";
		Trees_din <= x"009a1635";
		wait for Clk_period;
		Addr <=  "00010101110111";
		Trees_din <= x"ffb81635";
		wait for Clk_period;
		Addr <=  "00010101111000";
		Trees_din <= x"ffc01635";
		wait for Clk_period;
		Addr <=  "00010101111001";
		Trees_din <= x"0200f808";
		wait for Clk_period;
		Addr <=  "00010101111010";
		Trees_din <= x"1c002e04";
		wait for Clk_period;
		Addr <=  "00010101111011";
		Trees_din <= x"00d81635";
		wait for Clk_period;
		Addr <=  "00010101111100";
		Trees_din <= x"fff51635";
		wait for Clk_period;
		Addr <=  "00010101111101";
		Trees_din <= x"1b004208";
		wait for Clk_period;
		Addr <=  "00010101111110";
		Trees_din <= x"1b003604";
		wait for Clk_period;
		Addr <=  "00010101111111";
		Trees_din <= x"000f1635";
		wait for Clk_period;
		Addr <=  "00010110000000";
		Trees_din <= x"ffe21635";
		wait for Clk_period;
		Addr <=  "00010110000001";
		Trees_din <= x"11ff5404";
		wait for Clk_period;
		Addr <=  "00010110000010";
		Trees_din <= x"ffa11635";
		wait for Clk_period;
		Addr <=  "00010110000011";
		Trees_din <= x"00341635";
		wait for Clk_period;
		Addr <=  "00010110000100";
		Trees_din <= x"01076008";
		wait for Clk_period;
		Addr <=  "00010110000101";
		Trees_din <= x"02079804";
		wait for Clk_period;
		Addr <=  "00010110000110";
		Trees_din <= x"ff8e1635";
		wait for Clk_period;
		Addr <=  "00010110000111";
		Trees_din <= x"00281635";
		wait for Clk_period;
		Addr <=  "00010110001000";
		Trees_din <= x"03f86808";
		wait for Clk_period;
		Addr <=  "00010110001001";
		Trees_din <= x"07005104";
		wait for Clk_period;
		Addr <=  "00010110001010";
		Trees_din <= x"00661635";
		wait for Clk_period;
		Addr <=  "00010110001011";
		Trees_din <= x"ffb01635";
		wait for Clk_period;
		Addr <=  "00010110001100";
		Trees_din <= x"00ef1635";
		wait for Clk_period;
		Addr <=  "00010110001101";
		Trees_din <= x"11fab304";
		wait for Clk_period;
		Addr <=  "00010110001110";
		Trees_din <= x"ff8416f9";
		wait for Clk_period;
		Addr <=  "00010110001111";
		Trees_din <= x"02026c24";
		wait for Clk_period;
		Addr <=  "00010110010000";
		Trees_din <= x"03f89804";
		wait for Clk_period;
		Addr <=  "00010110010001";
		Trees_din <= x"ff7a16f9";
		wait for Clk_period;
		Addr <=  "00010110010010";
		Trees_din <= x"10056610";
		wait for Clk_period;
		Addr <=  "00010110010011";
		Trees_din <= x"13016808";
		wait for Clk_period;
		Addr <=  "00010110010100";
		Trees_din <= x"1d004704";
		wait for Clk_period;
		Addr <=  "00010110010101";
		Trees_din <= x"fff316f9";
		wait for Clk_period;
		Addr <=  "00010110010110";
		Trees_din <= x"ff8716f9";
		wait for Clk_period;
		Addr <=  "00010110010111";
		Trees_din <= x"10fb0804";
		wait for Clk_period;
		Addr <=  "00010110011000";
		Trees_din <= x"ffc516f9";
		wait for Clk_period;
		Addr <=  "00010110011001";
		Trees_din <= x"007e16f9";
		wait for Clk_period;
		Addr <=  "00010110011010";
		Trees_din <= x"0800ba08";
		wait for Clk_period;
		Addr <=  "00010110011011";
		Trees_din <= x"05fb6004";
		wait for Clk_period;
		Addr <=  "00010110011100";
		Trees_din <= x"000216f9";
		wait for Clk_period;
		Addr <=  "00010110011101";
		Trees_din <= x"00b016f9";
		wait for Clk_period;
		Addr <=  "00010110011110";
		Trees_din <= x"12fd9004";
		wait for Clk_period;
		Addr <=  "00010110011111";
		Trees_din <= x"008016f9";
		wait for Clk_period;
		Addr <=  "00010110100000";
		Trees_din <= x"ff8716f9";
		wait for Clk_period;
		Addr <=  "00010110100001";
		Trees_din <= x"00fe7b1c";
		wait for Clk_period;
		Addr <=  "00010110100010";
		Trees_din <= x"19009f0c";
		wait for Clk_period;
		Addr <=  "00010110100011";
		Trees_din <= x"13f86704";
		wait for Clk_period;
		Addr <=  "00010110100100";
		Trees_din <= x"ffa216f9";
		wait for Clk_period;
		Addr <=  "00010110100101";
		Trees_din <= x"0202d904";
		wait for Clk_period;
		Addr <=  "00010110100110";
		Trees_din <= x"ff9f16f9";
		wait for Clk_period;
		Addr <=  "00010110100111";
		Trees_din <= x"007c16f9";
		wait for Clk_period;
		Addr <=  "00010110101000";
		Trees_din <= x"1900a708";
		wait for Clk_period;
		Addr <=  "00010110101001";
		Trees_din <= x"0d010d04";
		wait for Clk_period;
		Addr <=  "00010110101010";
		Trees_din <= x"ffe216f9";
		wait for Clk_period;
		Addr <=  "00010110101011";
		Trees_din <= x"ff6c16f9";
		wait for Clk_period;
		Addr <=  "00010110101100";
		Trees_din <= x"10051404";
		wait for Clk_period;
		Addr <=  "00010110101101";
		Trees_din <= x"008416f9";
		wait for Clk_period;
		Addr <=  "00010110101110";
		Trees_din <= x"ffaf16f9";
		wait for Clk_period;
		Addr <=  "00010110101111";
		Trees_din <= x"0bf9f610";
		wait for Clk_period;
		Addr <=  "00010110110000";
		Trees_din <= x"0f00b308";
		wait for Clk_period;
		Addr <=  "00010110110001";
		Trees_din <= x"08022f04";
		wait for Clk_period;
		Addr <=  "00010110110010";
		Trees_din <= x"fffb16f9";
		wait for Clk_period;
		Addr <=  "00010110110011";
		Trees_din <= x"00a816f9";
		wait for Clk_period;
		Addr <=  "00010110110100";
		Trees_din <= x"0e020804";
		wait for Clk_period;
		Addr <=  "00010110110101";
		Trees_din <= x"ffee16f9";
		wait for Clk_period;
		Addr <=  "00010110110110";
		Trees_din <= x"ff6116f9";
		wait for Clk_period;
		Addr <=  "00010110110111";
		Trees_din <= x"1400ef08";
		wait for Clk_period;
		Addr <=  "00010110111000";
		Trees_din <= x"1400bb04";
		wait for Clk_period;
		Addr <=  "00010110111001";
		Trees_din <= x"000516f9";
		wait for Clk_period;
		Addr <=  "00010110111010";
		Trees_din <= x"ffa416f9";
		wait for Clk_period;
		Addr <=  "00010110111011";
		Trees_din <= x"16036304";
		wait for Clk_period;
		Addr <=  "00010110111100";
		Trees_din <= x"001316f9";
		wait for Clk_period;
		Addr <=  "00010110111101";
		Trees_din <= x"006b16f9";
		wait for Clk_period;
		Addr <=  "00010110111110";
		Trees_din <= x"0a03a348";
		wait for Clk_period;
		Addr <=  "00010110111111";
		Trees_din <= x"1104aa3c";
		wait for Clk_period;
		Addr <=  "00010111000000";
		Trees_din <= x"11043820";
		wait for Clk_period;
		Addr <=  "00010111000001";
		Trees_din <= x"0e025210";
		wait for Clk_period;
		Addr <=  "00010111000010";
		Trees_din <= x"1500ab08";
		wait for Clk_period;
		Addr <=  "00010111000011";
		Trees_din <= x"07005e04";
		wait for Clk_period;
		Addr <=  "00010111000100";
		Trees_din <= x"000b17ed";
		wait for Clk_period;
		Addr <=  "00010111000101";
		Trees_din <= x"ff8217ed";
		wait for Clk_period;
		Addr <=  "00010111000110";
		Trees_din <= x"14012e04";
		wait for Clk_period;
		Addr <=  "00010111000111";
		Trees_din <= x"008717ed";
		wait for Clk_period;
		Addr <=  "00010111001000";
		Trees_din <= x"ffd817ed";
		wait for Clk_period;
		Addr <=  "00010111001001";
		Trees_din <= x"0003e508";
		wait for Clk_period;
		Addr <=  "00010111001010";
		Trees_din <= x"07005704";
		wait for Clk_period;
		Addr <=  "00010111001011";
		Trees_din <= x"ffd317ed";
		wait for Clk_period;
		Addr <=  "00010111001100";
		Trees_din <= x"005c17ed";
		wait for Clk_period;
		Addr <=  "00010111001101";
		Trees_din <= x"0f007904";
		wait for Clk_period;
		Addr <=  "00010111001110";
		Trees_din <= x"001917ed";
		wait for Clk_period;
		Addr <=  "00010111001111";
		Trees_din <= x"ff8c17ed";
		wait for Clk_period;
		Addr <=  "00010111010000";
		Trees_din <= x"06f3df0c";
		wait for Clk_period;
		Addr <=  "00010111010001";
		Trees_din <= x"16003b04";
		wait for Clk_period;
		Addr <=  "00010111010010";
		Trees_din <= x"007f17ed";
		wait for Clk_period;
		Addr <=  "00010111010011";
		Trees_din <= x"0800d204";
		wait for Clk_period;
		Addr <=  "00010111010100";
		Trees_din <= x"ffdc17ed";
		wait for Clk_period;
		Addr <=  "00010111010101";
		Trees_din <= x"ff5b17ed";
		wait for Clk_period;
		Addr <=  "00010111010110";
		Trees_din <= x"02047508";
		wait for Clk_period;
		Addr <=  "00010111010111";
		Trees_din <= x"01049604";
		wait for Clk_period;
		Addr <=  "00010111011000";
		Trees_din <= x"004f17ed";
		wait for Clk_period;
		Addr <=  "00010111011001";
		Trees_din <= x"ff8e17ed";
		wait for Clk_period;
		Addr <=  "00010111011010";
		Trees_din <= x"09005404";
		wait for Clk_period;
		Addr <=  "00010111011011";
		Trees_din <= x"00ef17ed";
		wait for Clk_period;
		Addr <=  "00010111011100";
		Trees_din <= x"002a17ed";
		wait for Clk_period;
		Addr <=  "00010111011101";
		Trees_din <= x"020cbe08";
		wait for Clk_period;
		Addr <=  "00010111011110";
		Trees_din <= x"0afd2a04";
		wait for Clk_period;
		Addr <=  "00010111011111";
		Trees_din <= x"ff6817ed";
		wait for Clk_period;
		Addr <=  "00010111100000";
		Trees_din <= x"000417ed";
		wait for Clk_period;
		Addr <=  "00010111100001";
		Trees_din <= x"003d17ed";
		wait for Clk_period;
		Addr <=  "00010111100010";
		Trees_din <= x"0bf9f610";
		wait for Clk_period;
		Addr <=  "00010111100011";
		Trees_din <= x"03fda808";
		wait for Clk_period;
		Addr <=  "00010111100100";
		Trees_din <= x"1b003504";
		wait for Clk_period;
		Addr <=  "00010111100101";
		Trees_din <= x"ffdb17ed";
		wait for Clk_period;
		Addr <=  "00010111100110";
		Trees_din <= x"fee617ed";
		wait for Clk_period;
		Addr <=  "00010111100111";
		Trees_din <= x"16029b04";
		wait for Clk_period;
		Addr <=  "00010111101000";
		Trees_din <= x"ffbd17ed";
		wait for Clk_period;
		Addr <=  "00010111101001";
		Trees_din <= x"005217ed";
		wait for Clk_period;
		Addr <=  "00010111101010";
		Trees_din <= x"0e02b01c";
		wait for Clk_period;
		Addr <=  "00010111101011";
		Trees_din <= x"000ae810";
		wait for Clk_period;
		Addr <=  "00010111101100";
		Trees_din <= x"02068508";
		wait for Clk_period;
		Addr <=  "00010111101101";
		Trees_din <= x"05fdec04";
		wait for Clk_period;
		Addr <=  "00010111101110";
		Trees_din <= x"ff8d17ed";
		wait for Clk_period;
		Addr <=  "00010111101111";
		Trees_din <= x"007517ed";
		wait for Clk_period;
		Addr <=  "00010111110000";
		Trees_din <= x"0efe8604";
		wait for Clk_period;
		Addr <=  "00010111110001";
		Trees_din <= x"fffa17ed";
		wait for Clk_period;
		Addr <=  "00010111110010";
		Trees_din <= x"009417ed";
		wait for Clk_period;
		Addr <=  "00010111110011";
		Trees_din <= x"16003b04";
		wait for Clk_period;
		Addr <=  "00010111110100";
		Trees_din <= x"003117ed";
		wait for Clk_period;
		Addr <=  "00010111110101";
		Trees_din <= x"1500a504";
		wait for Clk_period;
		Addr <=  "00010111110110";
		Trees_din <= x"ff5117ed";
		wait for Clk_period;
		Addr <=  "00010111110111";
		Trees_din <= x"001a17ed";
		wait for Clk_period;
		Addr <=  "00010111111000";
		Trees_din <= x"1401b104";
		wait for Clk_period;
		Addr <=  "00010111111001";
		Trees_din <= x"00aa17ed";
		wait for Clk_period;
		Addr <=  "00010111111010";
		Trees_din <= x"001717ed";
		wait for Clk_period;
		Addr <=  "00010111111011";
		Trees_din <= x"02fce404";
		wait for Clk_period;
		Addr <=  "00010111111100";
		Trees_din <= x"ff8c1879";
		wait for Clk_period;
		Addr <=  "00010111111101";
		Trees_din <= x"11fab304";
		wait for Clk_period;
		Addr <=  "00010111111110";
		Trees_din <= x"ff8e1879";
		wait for Clk_period;
		Addr <=  "00010111111111";
		Trees_din <= x"1a00ac20";
		wait for Clk_period;
		Addr <=  "00011000000000";
		Trees_din <= x"1d004f10";
		wait for Clk_period;
		Addr <=  "00011000000001";
		Trees_din <= x"1c004708";
		wait for Clk_period;
		Addr <=  "00011000000010";
		Trees_din <= x"05f91a04";
		wait for Clk_period;
		Addr <=  "00011000000011";
		Trees_din <= x"ffaa1879";
		wait for Clk_period;
		Addr <=  "00011000000100";
		Trees_din <= x"005b1879";
		wait for Clk_period;
		Addr <=  "00011000000101";
		Trees_din <= x"0008bf04";
		wait for Clk_period;
		Addr <=  "00011000000110";
		Trees_din <= x"00331879";
		wait for Clk_period;
		Addr <=  "00011000000111";
		Trees_din <= x"01601879";
		wait for Clk_period;
		Addr <=  "00011000001000";
		Trees_din <= x"0f038408";
		wait for Clk_period;
		Addr <=  "00011000001001";
		Trees_din <= x"0b044904";
		wait for Clk_period;
		Addr <=  "00011000001010";
		Trees_din <= x"00391879";
		wait for Clk_period;
		Addr <=  "00011000001011";
		Trees_din <= x"ffb21879";
		wait for Clk_period;
		Addr <=  "00011000001100";
		Trees_din <= x"0c007a04";
		wait for Clk_period;
		Addr <=  "00011000001101";
		Trees_din <= x"fff31879";
		wait for Clk_period;
		Addr <=  "00011000001110";
		Trees_din <= x"ff5b1879";
		wait for Clk_period;
		Addr <=  "00011000001111";
		Trees_din <= x"18004510";
		wait for Clk_period;
		Addr <=  "00011000010000";
		Trees_din <= x"15008d08";
		wait for Clk_period;
		Addr <=  "00011000010001";
		Trees_din <= x"0efd4b04";
		wait for Clk_period;
		Addr <=  "00011000010010";
		Trees_din <= x"fff41879";
		wait for Clk_period;
		Addr <=  "00011000010011";
		Trees_din <= x"00a41879";
		wait for Clk_period;
		Addr <=  "00011000010100";
		Trees_din <= x"0110bb04";
		wait for Clk_period;
		Addr <=  "00011000010101";
		Trees_din <= x"00091879";
		wait for Clk_period;
		Addr <=  "00011000010110";
		Trees_din <= x"ffab1879";
		wait for Clk_period;
		Addr <=  "00011000010111";
		Trees_din <= x"03000c08";
		wait for Clk_period;
		Addr <=  "00011000011000";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00011000011001";
		Trees_din <= x"00201879";
		wait for Clk_period;
		Addr <=  "00011000011010";
		Trees_din <= x"ff8d1879";
		wait for Clk_period;
		Addr <=  "00011000011011";
		Trees_din <= x"1600db04";
		wait for Clk_period;
		Addr <=  "00011000011100";
		Trees_din <= x"ffef1879";
		wait for Clk_period;
		Addr <=  "00011000011101";
		Trees_din <= x"ff4e1879";
		wait for Clk_period;
		Addr <=  "00011000011110";
		Trees_din <= x"21000160";
		wait for Clk_period;
		Addr <=  "00011000011111";
		Trees_din <= x"1b002e28";
		wait for Clk_period;
		Addr <=  "00011000100000";
		Trees_din <= x"07005620";
		wait for Clk_period;
		Addr <=  "00011000100001";
		Trees_din <= x"02094410";
		wait for Clk_period;
		Addr <=  "00011000100010";
		Trees_din <= x"00097408";
		wait for Clk_period;
		Addr <=  "00011000100011";
		Trees_din <= x"08011d04";
		wait for Clk_period;
		Addr <=  "00011000100100";
		Trees_din <= x"00571965";
		wait for Clk_period;
		Addr <=  "00011000100101";
		Trees_din <= x"ffc21965";
		wait for Clk_period;
		Addr <=  "00011000100110";
		Trees_din <= x"16009f04";
		wait for Clk_period;
		Addr <=  "00011000100111";
		Trees_din <= x"ffe31965";
		wait for Clk_period;
		Addr <=  "00011000101000";
		Trees_din <= x"ff691965";
		wait for Clk_period;
		Addr <=  "00011000101001";
		Trees_din <= x"0d01f208";
		wait for Clk_period;
		Addr <=  "00011000101010";
		Trees_din <= x"0d00dd04";
		wait for Clk_period;
		Addr <=  "00011000101011";
		Trees_din <= x"00511965";
		wait for Clk_period;
		Addr <=  "00011000101100";
		Trees_din <= x"ffa61965";
		wait for Clk_period;
		Addr <=  "00011000101101";
		Trees_din <= x"1a00ff04";
		wait for Clk_period;
		Addr <=  "00011000101110";
		Trees_din <= x"00a21965";
		wait for Clk_period;
		Addr <=  "00011000101111";
		Trees_din <= x"000f1965";
		wait for Clk_period;
		Addr <=  "00011000110000";
		Trees_din <= x"07005804";
		wait for Clk_period;
		Addr <=  "00011000110001";
		Trees_din <= x"ff471965";
		wait for Clk_period;
		Addr <=  "00011000110010";
		Trees_din <= x"00391965";
		wait for Clk_period;
		Addr <=  "00011000110011";
		Trees_din <= x"1e006018";
		wait for Clk_period;
		Addr <=  "00011000110100";
		Trees_din <= x"08000908";
		wait for Clk_period;
		Addr <=  "00011000110101";
		Trees_din <= x"1b003104";
		wait for Clk_period;
		Addr <=  "00011000110110";
		Trees_din <= x"ff651965";
		wait for Clk_period;
		Addr <=  "00011000110111";
		Trees_din <= x"ffda1965";
		wait for Clk_period;
		Addr <=  "00011000111000";
		Trees_din <= x"0d002708";
		wait for Clk_period;
		Addr <=  "00011000111001";
		Trees_din <= x"06f36504";
		wait for Clk_period;
		Addr <=  "00011000111010";
		Trees_din <= x"ffe61965";
		wait for Clk_period;
		Addr <=  "00011000111011";
		Trees_din <= x"ff771965";
		wait for Clk_period;
		Addr <=  "00011000111100";
		Trees_din <= x"0b05a504";
		wait for Clk_period;
		Addr <=  "00011000111101";
		Trees_din <= x"004b1965";
		wait for Clk_period;
		Addr <=  "00011000111110";
		Trees_din <= x"ff861965";
		wait for Clk_period;
		Addr <=  "00011000111111";
		Trees_din <= x"1500a510";
		wait for Clk_period;
		Addr <=  "00011001000000";
		Trees_din <= x"1e006c08";
		wait for Clk_period;
		Addr <=  "00011001000001";
		Trees_din <= x"0800aa04";
		wait for Clk_period;
		Addr <=  "00011001000010";
		Trees_din <= x"ffa51965";
		wait for Clk_period;
		Addr <=  "00011001000011";
		Trees_din <= x"fff21965";
		wait for Clk_period;
		Addr <=  "00011001000100";
		Trees_din <= x"1e006d04";
		wait for Clk_period;
		Addr <=  "00011001000101";
		Trees_din <= x"00851965";
		wait for Clk_period;
		Addr <=  "00011001000110";
		Trees_din <= x"00001965";
		wait for Clk_period;
		Addr <=  "00011001000111";
		Trees_din <= x"1d003c08";
		wait for Clk_period;
		Addr <=  "00011001001000";
		Trees_din <= x"0c007104";
		wait for Clk_period;
		Addr <=  "00011001001001";
		Trees_din <= x"00401965";
		wait for Clk_period;
		Addr <=  "00011001001010";
		Trees_din <= x"ff931965";
		wait for Clk_period;
		Addr <=  "00011001001011";
		Trees_din <= x"0f003004";
		wait for Clk_period;
		Addr <=  "00011001001100";
		Trees_din <= x"001d1965";
		wait for Clk_period;
		Addr <=  "00011001001101";
		Trees_din <= x"00be1965";
		wait for Clk_period;
		Addr <=  "00011001001110";
		Trees_din <= x"01076008";
		wait for Clk_period;
		Addr <=  "00011001001111";
		Trees_din <= x"02079804";
		wait for Clk_period;
		Addr <=  "00011001010000";
		Trees_din <= x"ff8f1965";
		wait for Clk_period;
		Addr <=  "00011001010001";
		Trees_din <= x"00241965";
		wait for Clk_period;
		Addr <=  "00011001010010";
		Trees_din <= x"03f86808";
		wait for Clk_period;
		Addr <=  "00011001010011";
		Trees_din <= x"1c002904";
		wait for Clk_period;
		Addr <=  "00011001010100";
		Trees_din <= x"00641965";
		wait for Clk_period;
		Addr <=  "00011001010101";
		Trees_din <= x"ffb51965";
		wait for Clk_period;
		Addr <=  "00011001010110";
		Trees_din <= x"0afe5a04";
		wait for Clk_period;
		Addr <=  "00011001010111";
		Trees_din <= x"00d71965";
		wait for Clk_period;
		Addr <=  "00011001011000";
		Trees_din <= x"001c1965";
		wait for Clk_period;
		Addr <=  "00011001011001";
		Trees_din <= x"02047530";
		wait for Clk_period;
		Addr <=  "00011001011010";
		Trees_din <= x"03f89808";
		wait for Clk_period;
		Addr <=  "00011001011011";
		Trees_din <= x"1f000104";
		wait for Clk_period;
		Addr <=  "00011001011100";
		Trees_din <= x"ff761aa1";
		wait for Clk_period;
		Addr <=  "00011001011101";
		Trees_din <= x"00341aa1";
		wait for Clk_period;
		Addr <=  "00011001011110";
		Trees_din <= x"0ef96e0c";
		wait for Clk_period;
		Addr <=  "00011001011111";
		Trees_din <= x"1900a108";
		wait for Clk_period;
		Addr <=  "00011001100000";
		Trees_din <= x"05fcbb04";
		wait for Clk_period;
		Addr <=  "00011001100001";
		Trees_din <= x"ffa51aa1";
		wait for Clk_period;
		Addr <=  "00011001100010";
		Trees_din <= x"fff71aa1";
		wait for Clk_period;
		Addr <=  "00011001100011";
		Trees_din <= x"00f01aa1";
		wait for Clk_period;
		Addr <=  "00011001100100";
		Trees_din <= x"21000010";
		wait for Clk_period;
		Addr <=  "00011001100101";
		Trees_din <= x"03fd8408";
		wait for Clk_period;
		Addr <=  "00011001100110";
		Trees_din <= x"13f8d304";
		wait for Clk_period;
		Addr <=  "00011001100111";
		Trees_din <= x"00671aa1";
		wait for Clk_period;
		Addr <=  "00011001101000";
		Trees_din <= x"ff941aa1";
		wait for Clk_period;
		Addr <=  "00011001101001";
		Trees_din <= x"0e009f04";
		wait for Clk_period;
		Addr <=  "00011001101010";
		Trees_din <= x"ffce1aa1";
		wait for Clk_period;
		Addr <=  "00011001101011";
		Trees_din <= x"00161aa1";
		wait for Clk_period;
		Addr <=  "00011001101100";
		Trees_din <= x"15009204";
		wait for Clk_period;
		Addr <=  "00011001101101";
		Trees_din <= x"ff9f1aa1";
		wait for Clk_period;
		Addr <=  "00011001101110";
		Trees_din <= x"11005c04";
		wait for Clk_period;
		Addr <=  "00011001101111";
		Trees_din <= x"ffac1aa1";
		wait for Clk_period;
		Addr <=  "00011001110000";
		Trees_din <= x"00931aa1";
		wait for Clk_period;
		Addr <=  "00011001110001";
		Trees_din <= x"0802a538";
		wait for Clk_period;
		Addr <=  "00011001110010";
		Trees_din <= x"08020d1c";
		wait for Clk_period;
		Addr <=  "00011001110011";
		Trees_din <= x"0801b810";
		wait for Clk_period;
		Addr <=  "00011001110100";
		Trees_din <= x"11043808";
		wait for Clk_period;
		Addr <=  "00011001110101";
		Trees_din <= x"0e025a04";
		wait for Clk_period;
		Addr <=  "00011001110110";
		Trees_din <= x"00131aa1";
		wait for Clk_period;
		Addr <=  "00011001110111";
		Trees_din <= x"ffd21aa1";
		wait for Clk_period;
		Addr <=  "00011001111000";
		Trees_din <= x"09005404";
		wait for Clk_period;
		Addr <=  "00011001111001";
		Trees_din <= x"00a41aa1";
		wait for Clk_period;
		Addr <=  "00011001111010";
		Trees_din <= x"00021aa1";
		wait for Clk_period;
		Addr <=  "00011001111011";
		Trees_din <= x"10f74804";
		wait for Clk_period;
		Addr <=  "00011001111100";
		Trees_din <= x"00591aa1";
		wait for Clk_period;
		Addr <=  "00011001111101";
		Trees_din <= x"0afbee04";
		wait for Clk_period;
		Addr <=  "00011001111110";
		Trees_din <= x"000b1aa1";
		wait for Clk_period;
		Addr <=  "00011001111111";
		Trees_din <= x"ff801aa1";
		wait for Clk_period;
		Addr <=  "00011010000000";
		Trees_din <= x"11028410";
		wait for Clk_period;
		Addr <=  "00011010000001";
		Trees_din <= x"0206e308";
		wait for Clk_period;
		Addr <=  "00011010000010";
		Trees_din <= x"0a028404";
		wait for Clk_period;
		Addr <=  "00011010000011";
		Trees_din <= x"ff7b1aa1";
		wait for Clk_period;
		Addr <=  "00011010000100";
		Trees_din <= x"00151aa1";
		wait for Clk_period;
		Addr <=  "00011010000101";
		Trees_din <= x"1d004304";
		wait for Clk_period;
		Addr <=  "00011010000110";
		Trees_din <= x"009d1aa1";
		wait for Clk_period;
		Addr <=  "00011010000111";
		Trees_din <= x"fff11aa1";
		wait for Clk_period;
		Addr <=  "00011010001000";
		Trees_din <= x"08027708";
		wait for Clk_period;
		Addr <=  "00011010001001";
		Trees_din <= x"03f79304";
		wait for Clk_period;
		Addr <=  "00011010001010";
		Trees_din <= x"00371aa1";
		wait for Clk_period;
		Addr <=  "00011010001011";
		Trees_din <= x"00f51aa1";
		wait for Clk_period;
		Addr <=  "00011010001100";
		Trees_din <= x"00151aa1";
		wait for Clk_period;
		Addr <=  "00011010001101";
		Trees_din <= x"16027f1c";
		wait for Clk_period;
		Addr <=  "00011010001110";
		Trees_din <= x"10028710";
		wait for Clk_period;
		Addr <=  "00011010001111";
		Trees_din <= x"020abe08";
		wait for Clk_period;
		Addr <=  "00011010010000";
		Trees_din <= x"16025904";
		wait for Clk_period;
		Addr <=  "00011010010001";
		Trees_din <= x"ff701aa1";
		wait for Clk_period;
		Addr <=  "00011010010010";
		Trees_din <= x"00581aa1";
		wait for Clk_period;
		Addr <=  "00011010010011";
		Trees_din <= x"1c003304";
		wait for Clk_period;
		Addr <=  "00011010010100";
		Trees_din <= x"001a1aa1";
		wait for Clk_period;
		Addr <=  "00011010010101";
		Trees_din <= x"00751aa1";
		wait for Clk_period;
		Addr <=  "00011010010110";
		Trees_din <= x"0e00ab08";
		wait for Clk_period;
		Addr <=  "00011010010111";
		Trees_din <= x"09005304";
		wait for Clk_period;
		Addr <=  "00011010011000";
		Trees_din <= x"00251aa1";
		wait for Clk_period;
		Addr <=  "00011010011001";
		Trees_din <= x"00c51aa1";
		wait for Clk_period;
		Addr <=  "00011010011010";
		Trees_din <= x"fffa1aa1";
		wait for Clk_period;
		Addr <=  "00011010011011";
		Trees_din <= x"0700540c";
		wait for Clk_period;
		Addr <=  "00011010011100";
		Trees_din <= x"02080c04";
		wait for Clk_period;
		Addr <=  "00011010011101";
		Trees_din <= x"ff761aa1";
		wait for Clk_period;
		Addr <=  "00011010011110";
		Trees_din <= x"1e004b04";
		wait for Clk_period;
		Addr <=  "00011010011111";
		Trees_din <= x"ffb61aa1";
		wait for Clk_period;
		Addr <=  "00011010100000";
		Trees_din <= x"00691aa1";
		wait for Clk_period;
		Addr <=  "00011010100001";
		Trees_din <= x"0c020e08";
		wait for Clk_period;
		Addr <=  "00011010100010";
		Trees_din <= x"0d00a704";
		wait for Clk_period;
		Addr <=  "00011010100011";
		Trees_din <= x"ffdd1aa1";
		wait for Clk_period;
		Addr <=  "00011010100100";
		Trees_din <= x"ff2c1aa1";
		wait for Clk_period;
		Addr <=  "00011010100101";
		Trees_din <= x"1200a704";
		wait for Clk_period;
		Addr <=  "00011010100110";
		Trees_din <= x"00581aa1";
		wait for Clk_period;
		Addr <=  "00011010100111";
		Trees_din <= x"ff7d1aa1";
		wait for Clk_period;
		Addr <=  "00011010101000";
		Trees_din <= x"0406be6c";
		wait for Clk_period;
		Addr <=  "00011010101001";
		Trees_din <= x"0003e534";
		wait for Clk_period;
		Addr <=  "00011010101010";
		Trees_din <= x"010c4920";
		wait for Clk_period;
		Addr <=  "00011010101011";
		Trees_din <= x"05ff1810";
		wait for Clk_period;
		Addr <=  "00011010101100";
		Trees_din <= x"14020a08";
		wait for Clk_period;
		Addr <=  "00011010101101";
		Trees_din <= x"08022704";
		wait for Clk_period;
		Addr <=  "00011010101110";
		Trees_din <= x"00351bcd";
		wait for Clk_period;
		Addr <=  "00011010101111";
		Trees_din <= x"ffcf1bcd";
		wait for Clk_period;
		Addr <=  "00011010110000";
		Trees_din <= x"1b004604";
		wait for Clk_period;
		Addr <=  "00011010110001";
		Trees_din <= x"007b1bcd";
		wait for Clk_period;
		Addr <=  "00011010110010";
		Trees_din <= x"ffcd1bcd";
		wait for Clk_period;
		Addr <=  "00011010110011";
		Trees_din <= x"07005908";
		wait for Clk_period;
		Addr <=  "00011010110100";
		Trees_din <= x"0af7e104";
		wait for Clk_period;
		Addr <=  "00011010110101";
		Trees_din <= x"00441bcd";
		wait for Clk_period;
		Addr <=  "00011010110110";
		Trees_din <= x"ff7f1bcd";
		wait for Clk_period;
		Addr <=  "00011010110111";
		Trees_din <= x"0a017d04";
		wait for Clk_period;
		Addr <=  "00011010111000";
		Trees_din <= x"ffe11bcd";
		wait for Clk_period;
		Addr <=  "00011010111001";
		Trees_din <= x"00851bcd";
		wait for Clk_period;
		Addr <=  "00011010111010";
		Trees_din <= x"1900a50c";
		wait for Clk_period;
		Addr <=  "00011010111011";
		Trees_din <= x"00fae404";
		wait for Clk_period;
		Addr <=  "00011010111100";
		Trees_din <= x"002e1bcd";
		wait for Clk_period;
		Addr <=  "00011010111101";
		Trees_din <= x"0f000604";
		wait for Clk_period;
		Addr <=  "00011010111110";
		Trees_din <= x"ffdb1bcd";
		wait for Clk_period;
		Addr <=  "00011010111111";
		Trees_din <= x"ff681bcd";
		wait for Clk_period;
		Addr <=  "00011011000000";
		Trees_din <= x"1c002c04";
		wait for Clk_period;
		Addr <=  "00011011000001";
		Trees_din <= x"ffe11bcd";
		wait for Clk_period;
		Addr <=  "00011011000010";
		Trees_din <= x"00891bcd";
		wait for Clk_period;
		Addr <=  "00011011000011";
		Trees_din <= x"03fde01c";
		wait for Clk_period;
		Addr <=  "00011011000100";
		Trees_din <= x"06f0000c";
		wait for Clk_period;
		Addr <=  "00011011000101";
		Trees_din <= x"0009b104";
		wait for Clk_period;
		Addr <=  "00011011000110";
		Trees_din <= x"004d1bcd";
		wait for Clk_period;
		Addr <=  "00011011000111";
		Trees_din <= x"03f39604";
		wait for Clk_period;
		Addr <=  "00011011001000";
		Trees_din <= x"fffd1bcd";
		wait for Clk_period;
		Addr <=  "00011011001001";
		Trees_din <= x"ff5c1bcd";
		wait for Clk_period;
		Addr <=  "00011011001010";
		Trees_din <= x"0d032e08";
		wait for Clk_period;
		Addr <=  "00011011001011";
		Trees_din <= x"0d031204";
		wait for Clk_period;
		Addr <=  "00011011001100";
		Trees_din <= x"000d1bcd";
		wait for Clk_period;
		Addr <=  "00011011001101";
		Trees_din <= x"008c1bcd";
		wait for Clk_period;
		Addr <=  "00011011001110";
		Trees_din <= x"0f016804";
		wait for Clk_period;
		Addr <=  "00011011001111";
		Trees_din <= x"00091bcd";
		wait for Clk_period;
		Addr <=  "00011011010000";
		Trees_din <= x"ff7a1bcd";
		wait for Clk_period;
		Addr <=  "00011011010001";
		Trees_din <= x"1900820c";
		wait for Clk_period;
		Addr <=  "00011011010010";
		Trees_din <= x"03017908";
		wait for Clk_period;
		Addr <=  "00011011010011";
		Trees_din <= x"0d021404";
		wait for Clk_period;
		Addr <=  "00011011010100";
		Trees_din <= x"ffed1bcd";
		wait for Clk_period;
		Addr <=  "00011011010101";
		Trees_din <= x"00a71bcd";
		wait for Clk_period;
		Addr <=  "00011011010110";
		Trees_din <= x"ffa31bcd";
		wait for Clk_period;
		Addr <=  "00011011010111";
		Trees_din <= x"1e005508";
		wait for Clk_period;
		Addr <=  "00011011011000";
		Trees_din <= x"0201b304";
		wait for Clk_period;
		Addr <=  "00011011011001";
		Trees_din <= x"ff951bcd";
		wait for Clk_period;
		Addr <=  "00011011011010";
		Trees_din <= x"006e1bcd";
		wait for Clk_period;
		Addr <=  "00011011011011";
		Trees_din <= x"05fc3c04";
		wait for Clk_period;
		Addr <=  "00011011011100";
		Trees_din <= x"ffce1bcd";
		wait for Clk_period;
		Addr <=  "00011011011101";
		Trees_din <= x"ff591bcd";
		wait for Clk_period;
		Addr <=  "00011011011110";
		Trees_din <= x"0d032a1c";
		wait for Clk_period;
		Addr <=  "00011011011111";
		Trees_din <= x"1a00ac0c";
		wait for Clk_period;
		Addr <=  "00011011100000";
		Trees_din <= x"0f033b08";
		wait for Clk_period;
		Addr <=  "00011011100001";
		Trees_din <= x"00feee04";
		wait for Clk_period;
		Addr <=  "00011011100010";
		Trees_din <= x"ffed1bcd";
		wait for Clk_period;
		Addr <=  "00011011100011";
		Trees_din <= x"007d1bcd";
		wait for Clk_period;
		Addr <=  "00011011100100";
		Trees_din <= x"ffa81bcd";
		wait for Clk_period;
		Addr <=  "00011011100101";
		Trees_din <= x"1c002e04";
		wait for Clk_period;
		Addr <=  "00011011100110";
		Trees_din <= x"ff571bcd";
		wait for Clk_period;
		Addr <=  "00011011100111";
		Trees_din <= x"18004508";
		wait for Clk_period;
		Addr <=  "00011011101000";
		Trees_din <= x"17002904";
		wait for Clk_period;
		Addr <=  "00011011101001";
		Trees_din <= x"ffac1bcd";
		wait for Clk_period;
		Addr <=  "00011011101010";
		Trees_din <= x"003a1bcd";
		wait for Clk_period;
		Addr <=  "00011011101011";
		Trees_din <= x"ff6c1bcd";
		wait for Clk_period;
		Addr <=  "00011011101100";
		Trees_din <= x"07005704";
		wait for Clk_period;
		Addr <=  "00011011101101";
		Trees_din <= x"ffa61bcd";
		wait for Clk_period;
		Addr <=  "00011011101110";
		Trees_din <= x"14008004";
		wait for Clk_period;
		Addr <=  "00011011101111";
		Trees_din <= x"ffb91bcd";
		wait for Clk_period;
		Addr <=  "00011011110000";
		Trees_din <= x"1b003d04";
		wait for Clk_period;
		Addr <=  "00011011110001";
		Trees_din <= x"00c81bcd";
		wait for Clk_period;
		Addr <=  "00011011110010";
		Trees_din <= x"00291bcd";
		wait for Clk_period;
		Addr <=  "00011011110011";
		Trees_din <= x"0211fd6c";
		wait for Clk_period;
		Addr <=  "00011011110100";
		Trees_din <= x"1a00ac34";
		wait for Clk_period;
		Addr <=  "00011011110101";
		Trees_din <= x"1d004f1c";
		wait for Clk_period;
		Addr <=  "00011011110110";
		Trees_din <= x"06f40d0c";
		wait for Clk_period;
		Addr <=  "00011011110111";
		Trees_din <= x"0f03dc08";
		wait for Clk_period;
		Addr <=  "00011011111000";
		Trees_din <= x"08019304";
		wait for Clk_period;
		Addr <=  "00011011111001";
		Trees_din <= x"00c51cb9";
		wait for Clk_period;
		Addr <=  "00011011111010";
		Trees_din <= x"00121cb9";
		wait for Clk_period;
		Addr <=  "00011011111011";
		Trees_din <= x"ffb51cb9";
		wait for Clk_period;
		Addr <=  "00011011111100";
		Trees_din <= x"0c012008";
		wait for Clk_period;
		Addr <=  "00011011111101";
		Trees_din <= x"12006c04";
		wait for Clk_period;
		Addr <=  "00011011111110";
		Trees_din <= x"ffcf1cb9";
		wait for Clk_period;
		Addr <=  "00011011111111";
		Trees_din <= x"00a61cb9";
		wait for Clk_period;
		Addr <=  "00011100000000";
		Trees_din <= x"05fcdd04";
		wait for Clk_period;
		Addr <=  "00011100000001";
		Trees_din <= x"ff7d1cb9";
		wait for Clk_period;
		Addr <=  "00011100000010";
		Trees_din <= x"00321cb9";
		wait for Clk_period;
		Addr <=  "00011100000011";
		Trees_din <= x"0f038410";
		wait for Clk_period;
		Addr <=  "00011100000100";
		Trees_din <= x"08009108";
		wait for Clk_period;
		Addr <=  "00011100000101";
		Trees_din <= x"020d5c04";
		wait for Clk_period;
		Addr <=  "00011100000110";
		Trees_din <= x"ffd11cb9";
		wait for Clk_period;
		Addr <=  "00011100000111";
		Trees_din <= x"007d1cb9";
		wait for Clk_period;
		Addr <=  "00011100001000";
		Trees_din <= x"000e4f04";
		wait for Clk_period;
		Addr <=  "00011100001001";
		Trees_din <= x"00941cb9";
		wait for Clk_period;
		Addr <=  "00011100001010";
		Trees_din <= x"ffc31cb9";
		wait for Clk_period;
		Addr <=  "00011100001011";
		Trees_din <= x"0c007a04";
		wait for Clk_period;
		Addr <=  "00011100001100";
		Trees_din <= x"ffef1cb9";
		wait for Clk_period;
		Addr <=  "00011100001101";
		Trees_din <= x"ff631cb9";
		wait for Clk_period;
		Addr <=  "00011100001110";
		Trees_din <= x"1a00b618";
		wait for Clk_period;
		Addr <=  "00011100001111";
		Trees_din <= x"1401fb0c";
		wait for Clk_period;
		Addr <=  "00011100010000";
		Trees_din <= x"05fff708";
		wait for Clk_period;
		Addr <=  "00011100010001";
		Trees_din <= x"15008604";
		wait for Clk_period;
		Addr <=  "00011100010010";
		Trees_din <= x"ffea1cb9";
		wait for Clk_period;
		Addr <=  "00011100010011";
		Trees_din <= x"ff6b1cb9";
		wait for Clk_period;
		Addr <=  "00011100010100";
		Trees_din <= x"001a1cb9";
		wait for Clk_period;
		Addr <=  "00011100010101";
		Trees_din <= x"09005404";
		wait for Clk_period;
		Addr <=  "00011100010110";
		Trees_din <= x"ff691cb9";
		wait for Clk_period;
		Addr <=  "00011100010111";
		Trees_din <= x"14031004";
		wait for Clk_period;
		Addr <=  "00011100011000";
		Trees_din <= x"007c1cb9";
		wait for Clk_period;
		Addr <=  "00011100011001";
		Trees_din <= x"ffcf1cb9";
		wait for Clk_period;
		Addr <=  "00011100011010";
		Trees_din <= x"06f87f10";
		wait for Clk_period;
		Addr <=  "00011100011011";
		Trees_din <= x"0b04c108";
		wait for Clk_period;
		Addr <=  "00011100011100";
		Trees_din <= x"17006c04";
		wait for Clk_period;
		Addr <=  "00011100011101";
		Trees_din <= x"000a1cb9";
		wait for Clk_period;
		Addr <=  "00011100011110";
		Trees_din <= x"ffd31cb9";
		wait for Clk_period;
		Addr <=  "00011100011111";
		Trees_din <= x"0d027504";
		wait for Clk_period;
		Addr <=  "00011100100000";
		Trees_din <= x"00541cb9";
		wait for Clk_period;
		Addr <=  "00011100100001";
		Trees_din <= x"ffd91cb9";
		wait for Clk_period;
		Addr <=  "00011100100010";
		Trees_din <= x"18004108";
		wait for Clk_period;
		Addr <=  "00011100100011";
		Trees_din <= x"0d03a804";
		wait for Clk_period;
		Addr <=  "00011100100100";
		Trees_din <= x"00501cb9";
		wait for Clk_period;
		Addr <=  "00011100100101";
		Trees_din <= x"ff831cb9";
		wait for Clk_period;
		Addr <=  "00011100100110";
		Trees_din <= x"08002904";
		wait for Clk_period;
		Addr <=  "00011100100111";
		Trees_din <= x"00551cb9";
		wait for Clk_period;
		Addr <=  "00011100101000";
		Trees_din <= x"ffa71cb9";
		wait for Clk_period;
		Addr <=  "00011100101001";
		Trees_din <= x"17034f08";
		wait for Clk_period;
		Addr <=  "00011100101010";
		Trees_din <= x"0f039704";
		wait for Clk_period;
		Addr <=  "00011100101011";
		Trees_din <= x"00801cb9";
		wait for Clk_period;
		Addr <=  "00011100101100";
		Trees_din <= x"001f1cb9";
		wait for Clk_period;
		Addr <=  "00011100101101";
		Trees_din <= x"ffd01cb9";
		wait for Clk_period;
		Addr <=  "00011100101110";
		Trees_din <= x"02047538";
		wait for Clk_period;
		Addr <=  "00011100101111";
		Trees_din <= x"03f89808";
		wait for Clk_period;
		Addr <=  "00011100110000";
		Trees_din <= x"2003dd04";
		wait for Clk_period;
		Addr <=  "00011100110001";
		Trees_din <= x"00351dc5";
		wait for Clk_period;
		Addr <=  "00011100110010";
		Trees_din <= x"ff781dc5";
		wait for Clk_period;
		Addr <=  "00011100110011";
		Trees_din <= x"0ef96e10";
		wait for Clk_period;
		Addr <=  "00011100110100";
		Trees_din <= x"1900a108";
		wait for Clk_period;
		Addr <=  "00011100110101";
		Trees_din <= x"02004a04";
		wait for Clk_period;
		Addr <=  "00011100110110";
		Trees_din <= x"fff51dc5";
		wait for Clk_period;
		Addr <=  "00011100110111";
		Trees_din <= x"ffad1dc5";
		wait for Clk_period;
		Addr <=  "00011100111000";
		Trees_din <= x"1a00d704";
		wait for Clk_period;
		Addr <=  "00011100111001";
		Trees_din <= x"00ed1dc5";
		wait for Clk_period;
		Addr <=  "00011100111010";
		Trees_din <= x"00461dc5";
		wait for Clk_period;
		Addr <=  "00011100111011";
		Trees_din <= x"01fdfc10";
		wait for Clk_period;
		Addr <=  "00011100111100";
		Trees_din <= x"0c014c08";
		wait for Clk_period;
		Addr <=  "00011100111101";
		Trees_din <= x"01fb1904";
		wait for Clk_period;
		Addr <=  "00011100111110";
		Trees_din <= x"00741dc5";
		wait for Clk_period;
		Addr <=  "00011100111111";
		Trees_din <= x"ffb91dc5";
		wait for Clk_period;
		Addr <=  "00011101000000";
		Trees_din <= x"1301c404";
		wait for Clk_period;
		Addr <=  "00011101000001";
		Trees_din <= x"ff6f1dc5";
		wait for Clk_period;
		Addr <=  "00011101000010";
		Trees_din <= x"fffb1dc5";
		wait for Clk_period;
		Addr <=  "00011101000011";
		Trees_din <= x"16009408";
		wait for Clk_period;
		Addr <=  "00011101000100";
		Trees_din <= x"21000004";
		wait for Clk_period;
		Addr <=  "00011101000101";
		Trees_din <= x"ffa51dc5";
		wait for Clk_period;
		Addr <=  "00011101000110";
		Trees_din <= x"00431dc5";
		wait for Clk_period;
		Addr <=  "00011101000111";
		Trees_din <= x"1900a304";
		wait for Clk_period;
		Addr <=  "00011101001000";
		Trees_din <= x"00251dc5";
		wait for Clk_period;
		Addr <=  "00011101001001";
		Trees_din <= x"ffca1dc5";
		wait for Clk_period;
		Addr <=  "00011101001010";
		Trees_din <= x"0e041138";
		wait for Clk_period;
		Addr <=  "00011101001011";
		Trees_din <= x"11044420";
		wait for Clk_period;
		Addr <=  "00011101001100";
		Trees_din <= x"00fe7b10";
		wait for Clk_period;
		Addr <=  "00011101001101";
		Trees_din <= x"0e005a08";
		wait for Clk_period;
		Addr <=  "00011101001110";
		Trees_din <= x"07005b04";
		wait for Clk_period;
		Addr <=  "00011101001111";
		Trees_din <= x"ffcd1dc5";
		wait for Clk_period;
		Addr <=  "00011101010000";
		Trees_din <= x"00631dc5";
		wait for Clk_period;
		Addr <=  "00011101010001";
		Trees_din <= x"05f6a104";
		wait for Clk_period;
		Addr <=  "00011101010010";
		Trees_din <= x"000c1dc5";
		wait for Clk_period;
		Addr <=  "00011101010011";
		Trees_din <= x"00a31dc5";
		wait for Clk_period;
		Addr <=  "00011101010100";
		Trees_din <= x"0e025a08";
		wait for Clk_period;
		Addr <=  "00011101010101";
		Trees_din <= x"11030f04";
		wait for Clk_period;
		Addr <=  "00011101010110";
		Trees_din <= x"00081dc5";
		wait for Clk_period;
		Addr <=  "00011101010111";
		Trees_din <= x"00991dc5";
		wait for Clk_period;
		Addr <=  "00011101011000";
		Trees_din <= x"06f87f04";
		wait for Clk_period;
		Addr <=  "00011101011001";
		Trees_din <= x"ffb81dc5";
		wait for Clk_period;
		Addr <=  "00011101011010";
		Trees_din <= x"00551dc5";
		wait for Clk_period;
		Addr <=  "00011101011011";
		Trees_din <= x"06f4d30c";
		wait for Clk_period;
		Addr <=  "00011101011100";
		Trees_din <= x"1401dd08";
		wait for Clk_period;
		Addr <=  "00011101011101";
		Trees_din <= x"0c011904";
		wait for Clk_period;
		Addr <=  "00011101011110";
		Trees_din <= x"00101dc5";
		wait for Clk_period;
		Addr <=  "00011101011111";
		Trees_din <= x"ff8b1dc5";
		wait for Clk_period;
		Addr <=  "00011101100000";
		Trees_din <= x"00561dc5";
		wait for Clk_period;
		Addr <=  "00011101100001";
		Trees_din <= x"06fa9b08";
		wait for Clk_period;
		Addr <=  "00011101100010";
		Trees_din <= x"10facc04";
		wait for Clk_period;
		Addr <=  "00011101100011";
		Trees_din <= x"00251dc5";
		wait for Clk_period;
		Addr <=  "00011101100100";
		Trees_din <= x"00e11dc5";
		wait for Clk_period;
		Addr <=  "00011101100101";
		Trees_din <= x"ffdd1dc5";
		wait for Clk_period;
		Addr <=  "00011101100110";
		Trees_din <= x"10fade08";
		wait for Clk_period;
		Addr <=  "00011101100111";
		Trees_din <= x"0d01ce04";
		wait for Clk_period;
		Addr <=  "00011101101000";
		Trees_din <= x"00701dc5";
		wait for Clk_period;
		Addr <=  "00011101101001";
		Trees_din <= x"ffc81dc5";
		wait for Clk_period;
		Addr <=  "00011101101010";
		Trees_din <= x"0f007b04";
		wait for Clk_period;
		Addr <=  "00011101101011";
		Trees_din <= x"002f1dc5";
		wait for Clk_period;
		Addr <=  "00011101101100";
		Trees_din <= x"0f025f04";
		wait for Clk_period;
		Addr <=  "00011101101101";
		Trees_din <= x"ff551dc5";
		wait for Clk_period;
		Addr <=  "00011101101110";
		Trees_din <= x"14032404";
		wait for Clk_period;
		Addr <=  "00011101101111";
		Trees_din <= x"00311dc5";
		wait for Clk_period;
		Addr <=  "00011101110000";
		Trees_din <= x"ffa11dc5";
		wait for Clk_period;
		Addr <=  "00011101110001";
		Trees_din <= x"0a03a35c";
		wait for Clk_period;
		Addr <=  "00011101110010";
		Trees_din <= x"04f95834";
		wait for Clk_period;
		Addr <=  "00011101110011";
		Trees_din <= x"020baf1c";
		wait for Clk_period;
		Addr <=  "00011101110100";
		Trees_din <= x"1800380c";
		wait for Clk_period;
		Addr <=  "00011101110101";
		Trees_din <= x"1a00ef08";
		wait for Clk_period;
		Addr <=  "00011101110110";
		Trees_din <= x"010b3204";
		wait for Clk_period;
		Addr <=  "00011101110111";
		Trees_din <= x"001d1ee1";
		wait for Clk_period;
		Addr <=  "00011101111000";
		Trees_din <= x"00c01ee1";
		wait for Clk_period;
		Addr <=  "00011101111001";
		Trees_din <= x"ffb61ee1";
		wait for Clk_period;
		Addr <=  "00011101111010";
		Trees_din <= x"1c004008";
		wait for Clk_period;
		Addr <=  "00011101111011";
		Trees_din <= x"13015e04";
		wait for Clk_period;
		Addr <=  "00011101111100";
		Trees_din <= x"ff901ee1";
		wait for Clk_period;
		Addr <=  "00011101111101";
		Trees_din <= x"00231ee1";
		wait for Clk_period;
		Addr <=  "00011101111110";
		Trees_din <= x"1e008504";
		wait for Clk_period;
		Addr <=  "00011101111111";
		Trees_din <= x"00561ee1";
		wait for Clk_period;
		Addr <=  "00011110000000";
		Trees_din <= x"ffa71ee1";
		wait for Clk_period;
		Addr <=  "00011110000001";
		Trees_din <= x"0d032a0c";
		wait for Clk_period;
		Addr <=  "00011110000010";
		Trees_din <= x"0af77a04";
		wait for Clk_period;
		Addr <=  "00011110000011";
		Trees_din <= x"ff9f1ee1";
		wait for Clk_period;
		Addr <=  "00011110000100";
		Trees_din <= x"09005104";
		wait for Clk_period;
		Addr <=  "00011110000101";
		Trees_din <= x"000e1ee1";
		wait for Clk_period;
		Addr <=  "00011110000110";
		Trees_din <= x"00911ee1";
		wait for Clk_period;
		Addr <=  "00011110000111";
		Trees_din <= x"1401ad08";
		wait for Clk_period;
		Addr <=  "00011110001000";
		Trees_din <= x"16037804";
		wait for Clk_period;
		Addr <=  "00011110001001";
		Trees_din <= x"00691ee1";
		wait for Clk_period;
		Addr <=  "00011110001010";
		Trees_din <= x"ffa41ee1";
		wait for Clk_period;
		Addr <=  "00011110001011";
		Trees_din <= x"ff4a1ee1";
		wait for Clk_period;
		Addr <=  "00011110001100";
		Trees_din <= x"04f9a008";
		wait for Clk_period;
		Addr <=  "00011110001101";
		Trees_din <= x"0205dc04";
		wait for Clk_period;
		Addr <=  "00011110001110";
		Trees_din <= x"ffff1ee1";
		wait for Clk_period;
		Addr <=  "00011110001111";
		Trees_din <= x"00971ee1";
		wait for Clk_period;
		Addr <=  "00011110010000";
		Trees_din <= x"05fbe610";
		wait for Clk_period;
		Addr <=  "00011110010001";
		Trees_din <= x"15009e08";
		wait for Clk_period;
		Addr <=  "00011110010010";
		Trees_din <= x"02ff5f04";
		wait for Clk_period;
		Addr <=  "00011110010011";
		Trees_din <= x"ff8c1ee1";
		wait for Clk_period;
		Addr <=  "00011110010100";
		Trees_din <= x"003a1ee1";
		wait for Clk_period;
		Addr <=  "00011110010101";
		Trees_din <= x"03024704";
		wait for Clk_period;
		Addr <=  "00011110010110";
		Trees_din <= x"ffc41ee1";
		wait for Clk_period;
		Addr <=  "00011110010111";
		Trees_din <= x"003b1ee1";
		wait for Clk_period;
		Addr <=  "00011110011000";
		Trees_din <= x"04012008";
		wait for Clk_period;
		Addr <=  "00011110011001";
		Trees_din <= x"05fcc804";
		wait for Clk_period;
		Addr <=  "00011110011010";
		Trees_din <= x"ff8d1ee1";
		wait for Clk_period;
		Addr <=  "00011110011011";
		Trees_din <= x"fff51ee1";
		wait for Clk_period;
		Addr <=  "00011110011100";
		Trees_din <= x"0f008604";
		wait for Clk_period;
		Addr <=  "00011110011101";
		Trees_din <= x"ffdf1ee1";
		wait for Clk_period;
		Addr <=  "00011110011110";
		Trees_din <= x"00341ee1";
		wait for Clk_period;
		Addr <=  "00011110011111";
		Trees_din <= x"0bf9f610";
		wait for Clk_period;
		Addr <=  "00011110100000";
		Trees_din <= x"03fda808";
		wait for Clk_period;
		Addr <=  "00011110100001";
		Trees_din <= x"03f9d604";
		wait for Clk_period;
		Addr <=  "00011110100010";
		Trees_din <= x"ffd31ee1";
		wait for Clk_period;
		Addr <=  "00011110100011";
		Trees_din <= x"ff171ee1";
		wait for Clk_period;
		Addr <=  "00011110100100";
		Trees_din <= x"0d02a704";
		wait for Clk_period;
		Addr <=  "00011110100101";
		Trees_din <= x"002d1ee1";
		wait for Clk_period;
		Addr <=  "00011110100110";
		Trees_din <= x"ffce1ee1";
		wait for Clk_period;
		Addr <=  "00011110100111";
		Trees_din <= x"0e02b01c";
		wait for Clk_period;
		Addr <=  "00011110101000";
		Trees_din <= x"000ae810";
		wait for Clk_period;
		Addr <=  "00011110101001";
		Trees_din <= x"17000208";
		wait for Clk_period;
		Addr <=  "00011110101010";
		Trees_din <= x"0201c104";
		wait for Clk_period;
		Addr <=  "00011110101011";
		Trees_din <= x"ffd21ee1";
		wait for Clk_period;
		Addr <=  "00011110101100";
		Trees_din <= x"00751ee1";
		wait for Clk_period;
		Addr <=  "00011110101101";
		Trees_din <= x"02089504";
		wait for Clk_period;
		Addr <=  "00011110101110";
		Trees_din <= x"ff891ee1";
		wait for Clk_period;
		Addr <=  "00011110101111";
		Trees_din <= x"00611ee1";
		wait for Clk_period;
		Addr <=  "00011110110000";
		Trees_din <= x"1a00f108";
		wait for Clk_period;
		Addr <=  "00011110110001";
		Trees_din <= x"12fd7304";
		wait for Clk_period;
		Addr <=  "00011110110010";
		Trees_din <= x"00001ee1";
		wait for Clk_period;
		Addr <=  "00011110110011";
		Trees_din <= x"ff631ee1";
		wait for Clk_period;
		Addr <=  "00011110110100";
		Trees_din <= x"00501ee1";
		wait for Clk_period;
		Addr <=  "00011110110101";
		Trees_din <= x"02071404";
		wait for Clk_period;
		Addr <=  "00011110110110";
		Trees_din <= x"00231ee1";
		wait for Clk_period;
		Addr <=  "00011110110111";
		Trees_din <= x"00921ee1";
		wait for Clk_period;
		Addr <=  "00011110111000";
		Trees_din <= x"0208324c";
		wait for Clk_period;
		Addr <=  "00011110111001";
		Trees_din <= x"010f7440";
		wait for Clk_period;
		Addr <=  "00011110111010";
		Trees_din <= x"0d037b20";
		wait for Clk_period;
		Addr <=  "00011110111011";
		Trees_din <= x"08017510";
		wait for Clk_period;
		Addr <=  "00011110111100";
		Trees_din <= x"010d2808";
		wait for Clk_period;
		Addr <=  "00011110111101";
		Trees_din <= x"1d004604";
		wait for Clk_period;
		Addr <=  "00011110111110";
		Trees_din <= x"00281fd5";
		wait for Clk_period;
		Addr <=  "00011110111111";
		Trees_din <= x"ffe01fd5";
		wait for Clk_period;
		Addr <=  "00011111000000";
		Trees_din <= x"11027304";
		wait for Clk_period;
		Addr <=  "00011111000001";
		Trees_din <= x"00b71fd5";
		wait for Clk_period;
		Addr <=  "00011111000010";
		Trees_din <= x"ffda1fd5";
		wait for Clk_period;
		Addr <=  "00011111000011";
		Trees_din <= x"0801f408";
		wait for Clk_period;
		Addr <=  "00011111000100";
		Trees_din <= x"1603e104";
		wait for Clk_period;
		Addr <=  "00011111000101";
		Trees_din <= x"ff8e1fd5";
		wait for Clk_period;
		Addr <=  "00011111000110";
		Trees_din <= x"00281fd5";
		wait for Clk_period;
		Addr <=  "00011111000111";
		Trees_din <= x"0204f604";
		wait for Clk_period;
		Addr <=  "00011111001000";
		Trees_din <= x"00211fd5";
		wait for Clk_period;
		Addr <=  "00011111001001";
		Trees_din <= x"ffc61fd5";
		wait for Clk_period;
		Addr <=  "00011111001010";
		Trees_din <= x"07005710";
		wait for Clk_period;
		Addr <=  "00011111001011";
		Trees_din <= x"0f003f08";
		wait for Clk_period;
		Addr <=  "00011111001100";
		Trees_din <= x"14010d04";
		wait for Clk_period;
		Addr <=  "00011111001101";
		Trees_din <= x"ffb91fd5";
		wait for Clk_period;
		Addr <=  "00011111001110";
		Trees_din <= x"003f1fd5";
		wait for Clk_period;
		Addr <=  "00011111001111";
		Trees_din <= x"1a00a304";
		wait for Clk_period;
		Addr <=  "00011111010000";
		Trees_din <= x"ffd41fd5";
		wait for Clk_period;
		Addr <=  "00011111010001";
		Trees_din <= x"ff5e1fd5";
		wait for Clk_period;
		Addr <=  "00011111010010";
		Trees_din <= x"00046408";
		wait for Clk_period;
		Addr <=  "00011111010011";
		Trees_din <= x"0d03db04";
		wait for Clk_period;
		Addr <=  "00011111010100";
		Trees_din <= x"00771fd5";
		wait for Clk_period;
		Addr <=  "00011111010101";
		Trees_din <= x"ffd51fd5";
		wait for Clk_period;
		Addr <=  "00011111010110";
		Trees_din <= x"1203f704";
		wait for Clk_period;
		Addr <=  "00011111010111";
		Trees_din <= x"ff8a1fd5";
		wait for Clk_period;
		Addr <=  "00011111011000";
		Trees_din <= x"005e1fd5";
		wait for Clk_period;
		Addr <=  "00011111011001";
		Trees_din <= x"05fb6b08";
		wait for Clk_period;
		Addr <=  "00011111011010";
		Trees_din <= x"11046804";
		wait for Clk_period;
		Addr <=  "00011111011011";
		Trees_din <= x"ff711fd5";
		wait for Clk_period;
		Addr <=  "00011111011100";
		Trees_din <= x"00441fd5";
		wait for Clk_period;
		Addr <=  "00011111011101";
		Trees_din <= x"00591fd5";
		wait for Clk_period;
		Addr <=  "00011111011110";
		Trees_din <= x"0800050c";
		wait for Clk_period;
		Addr <=  "00011111011111";
		Trees_din <= x"07005908";
		wait for Clk_period;
		Addr <=  "00011111100000";
		Trees_din <= x"020b6104";
		wait for Clk_period;
		Addr <=  "00011111100001";
		Trees_din <= x"ffc01fd5";
		wait for Clk_period;
		Addr <=  "00011111100010";
		Trees_din <= x"00711fd5";
		wait for Clk_period;
		Addr <=  "00011111100011";
		Trees_din <= x"00951fd5";
		wait for Clk_period;
		Addr <=  "00011111100100";
		Trees_din <= x"1006831c";
		wait for Clk_period;
		Addr <=  "00011111100101";
		Trees_din <= x"04f6740c";
		wait for Clk_period;
		Addr <=  "00011111100110";
		Trees_din <= x"10f9dc04";
		wait for Clk_period;
		Addr <=  "00011111100111";
		Trees_din <= x"ffca1fd5";
		wait for Clk_period;
		Addr <=  "00011111101000";
		Trees_din <= x"10054e04";
		wait for Clk_period;
		Addr <=  "00011111101001";
		Trees_din <= x"00791fd5";
		wait for Clk_period;
		Addr <=  "00011111101010";
		Trees_din <= x"ffdd1fd5";
		wait for Clk_period;
		Addr <=  "00011111101011";
		Trees_din <= x"10f9a208";
		wait for Clk_period;
		Addr <=  "00011111101100";
		Trees_din <= x"010b7604";
		wait for Clk_period;
		Addr <=  "00011111101101";
		Trees_din <= x"00761fd5";
		wait for Clk_period;
		Addr <=  "00011111101110";
		Trees_din <= x"ffbf1fd5";
		wait for Clk_period;
		Addr <=  "00011111101111";
		Trees_din <= x"03fe8b04";
		wait for Clk_period;
		Addr <=  "00011111110000";
		Trees_din <= x"ffe51fd5";
		wait for Clk_period;
		Addr <=  "00011111110001";
		Trees_din <= x"003c1fd5";
		wait for Clk_period;
		Addr <=  "00011111110010";
		Trees_din <= x"01070104";
		wait for Clk_period;
		Addr <=  "00011111110011";
		Trees_din <= x"002c1fd5";
		wait for Clk_period;
		Addr <=  "00011111110100";
		Trees_din <= x"00941fd5";
		wait for Clk_period;
		Addr <=  "00011111110101";
		Trees_din <= x"0204752c";
		wait for Clk_period;
		Addr <=  "00011111110110";
		Trees_din <= x"03fa3610";
		wait for Clk_period;
		Addr <=  "00011111110111";
		Trees_din <= x"0b05670c";
		wait for Clk_period;
		Addr <=  "00011111111000";
		Trees_din <= x"12fd9004";
		wait for Clk_period;
		Addr <=  "00011111111001";
		Trees_din <= x"001320f9";
		wait for Clk_period;
		Addr <=  "00011111111010";
		Trees_din <= x"0006ac04";
		wait for Clk_period;
		Addr <=  "00011111111011";
		Trees_din <= x"fff720f9";
		wait for Clk_period;
		Addr <=  "00011111111100";
		Trees_din <= x"ff7720f9";
		wait for Clk_period;
		Addr <=  "00011111111101";
		Trees_din <= x"004b20f9";
		wait for Clk_period;
		Addr <=  "00011111111110";
		Trees_din <= x"0ef96e0c";
		wait for Clk_period;
		Addr <=  "00011111111111";
		Trees_din <= x"1900a104";
		wait for Clk_period;
		Addr <=  "00100000000000";
		Trees_din <= x"ffc220f9";
		wait for Clk_period;
		Addr <=  "00100000000001";
		Trees_din <= x"0c026804";
		wait for Clk_period;
		Addr <=  "00100000000010";
		Trees_din <= x"003520f9";
		wait for Clk_period;
		Addr <=  "00100000000011";
		Trees_din <= x"00d620f9";
		wait for Clk_period;
		Addr <=  "00100000000100";
		Trees_din <= x"000f360c";
		wait for Clk_period;
		Addr <=  "00100000000101";
		Trees_din <= x"000e9008";
		wait for Clk_period;
		Addr <=  "00100000000110";
		Trees_din <= x"1a00a204";
		wait for Clk_period;
		Addr <=  "00100000000111";
		Trees_din <= x"003220f9";
		wait for Clk_period;
		Addr <=  "00100000001000";
		Trees_din <= x"ffe820f9";
		wait for Clk_period;
		Addr <=  "00100000001001";
		Trees_din <= x"008a20f9";
		wait for Clk_period;
		Addr <=  "00100000001010";
		Trees_din <= x"ff8820f9";
		wait for Clk_period;
		Addr <=  "00100000001011";
		Trees_din <= x"13f92e2c";
		wait for Clk_period;
		Addr <=  "00100000001100";
		Trees_din <= x"19009e1c";
		wait for Clk_period;
		Addr <=  "00100000001101";
		Trees_din <= x"03f94d10";
		wait for Clk_period;
		Addr <=  "00100000001110";
		Trees_din <= x"13f88008";
		wait for Clk_period;
		Addr <=  "00100000001111";
		Trees_din <= x"05fca304";
		wait for Clk_period;
		Addr <=  "00100000010000";
		Trees_din <= x"000d20f9";
		wait for Clk_period;
		Addr <=  "00100000010001";
		Trees_din <= x"005120f9";
		wait for Clk_period;
		Addr <=  "00100000010010";
		Trees_din <= x"09005404";
		wait for Clk_period;
		Addr <=  "00100000010011";
		Trees_din <= x"ffe420f9";
		wait for Clk_period;
		Addr <=  "00100000010100";
		Trees_din <= x"ff6120f9";
		wait for Clk_period;
		Addr <=  "00100000010101";
		Trees_din <= x"13f86f04";
		wait for Clk_period;
		Addr <=  "00100000010110";
		Trees_din <= x"ffb620f9";
		wait for Clk_period;
		Addr <=  "00100000010111";
		Trees_din <= x"05faab04";
		wait for Clk_period;
		Addr <=  "00100000011000";
		Trees_din <= x"001820f9";
		wait for Clk_period;
		Addr <=  "00100000011001";
		Trees_din <= x"00a920f9";
		wait for Clk_period;
		Addr <=  "00100000011010";
		Trees_din <= x"18003704";
		wait for Clk_period;
		Addr <=  "00100000011011";
		Trees_din <= x"003120f9";
		wait for Clk_period;
		Addr <=  "00100000011100";
		Trees_din <= x"13f88904";
		wait for Clk_period;
		Addr <=  "00100000011101";
		Trees_din <= x"fffe20f9";
		wait for Clk_period;
		Addr <=  "00100000011110";
		Trees_din <= x"09004f04";
		wait for Clk_period;
		Addr <=  "00100000011111";
		Trees_din <= x"ffe720f9";
		wait for Clk_period;
		Addr <=  "00100000100000";
		Trees_din <= x"ff4f20f9";
		wait for Clk_period;
		Addr <=  "00100000100001";
		Trees_din <= x"12005e1c";
		wait for Clk_period;
		Addr <=  "00100000100010";
		Trees_din <= x"0800540c";
		wait for Clk_period;
		Addr <=  "00100000100011";
		Trees_din <= x"0e008f08";
		wait for Clk_period;
		Addr <=  "00100000100100";
		Trees_din <= x"0d019304";
		wait for Clk_period;
		Addr <=  "00100000100101";
		Trees_din <= x"fff720f9";
		wait for Clk_period;
		Addr <=  "00100000100110";
		Trees_din <= x"ff6320f9";
		wait for Clk_period;
		Addr <=  "00100000100111";
		Trees_din <= x"004b20f9";
		wait for Clk_period;
		Addr <=  "00100000101000";
		Trees_din <= x"0b034308";
		wait for Clk_period;
		Addr <=  "00100000101001";
		Trees_din <= x"12fef604";
		wait for Clk_period;
		Addr <=  "00100000101010";
		Trees_din <= x"ffd520f9";
		wait for Clk_period;
		Addr <=  "00100000101011";
		Trees_din <= x"004e20f9";
		wait for Clk_period;
		Addr <=  "00100000101100";
		Trees_din <= x"08011a04";
		wait for Clk_period;
		Addr <=  "00100000101101";
		Trees_din <= x"00b020f9";
		wait for Clk_period;
		Addr <=  "00100000101110";
		Trees_din <= x"002c20f9";
		wait for Clk_period;
		Addr <=  "00100000101111";
		Trees_din <= x"16003b10";
		wait for Clk_period;
		Addr <=  "00100000110000";
		Trees_din <= x"0c00d308";
		wait for Clk_period;
		Addr <=  "00100000110001";
		Trees_din <= x"0105bc04";
		wait for Clk_period;
		Addr <=  "00100000110010";
		Trees_din <= x"003d20f9";
		wait for Clk_period;
		Addr <=  "00100000110011";
		Trees_din <= x"ff8920f9";
		wait for Clk_period;
		Addr <=  "00100000110100";
		Trees_din <= x"15009d04";
		wait for Clk_period;
		Addr <=  "00100000110101";
		Trees_din <= x"007f20f9";
		wait for Clk_period;
		Addr <=  "00100000110110";
		Trees_din <= x"ffd220f9";
		wait for Clk_period;
		Addr <=  "00100000110111";
		Trees_din <= x"0c02c108";
		wait for Clk_period;
		Addr <=  "00100000111000";
		Trees_din <= x"11000d04";
		wait for Clk_period;
		Addr <=  "00100000111001";
		Trees_din <= x"ff8920f9";
		wait for Clk_period;
		Addr <=  "00100000111010";
		Trees_din <= x"001320f9";
		wait for Clk_period;
		Addr <=  "00100000111011";
		Trees_din <= x"19009404";
		wait for Clk_period;
		Addr <=  "00100000111100";
		Trees_din <= x"ffa020f9";
		wait for Clk_period;
		Addr <=  "00100000111101";
		Trees_din <= x"000420f9";
		wait for Clk_period;
		Addr <=  "00100000111110";
		Trees_din <= x"03f40e14";
		wait for Clk_period;
		Addr <=  "00100000111111";
		Trees_din <= x"020e8d0c";
		wait for Clk_period;
		Addr <=  "00100001000000";
		Trees_din <= x"09005a08";
		wait for Clk_period;
		Addr <=  "00100001000001";
		Trees_din <= x"1b003204";
		wait for Clk_period;
		Addr <=  "00100001000010";
		Trees_din <= x"ffe72185";
		wait for Clk_period;
		Addr <=  "00100001000011";
		Trees_din <= x"ff782185";
		wait for Clk_period;
		Addr <=  "00100001000100";
		Trees_din <= x"001c2185";
		wait for Clk_period;
		Addr <=  "00100001000101";
		Trees_din <= x"0bfa8104";
		wait for Clk_period;
		Addr <=  "00100001000110";
		Trees_din <= x"005c2185";
		wait for Clk_period;
		Addr <=  "00100001000111";
		Trees_din <= x"ffdf2185";
		wait for Clk_period;
		Addr <=  "00100001001000";
		Trees_din <= x"03f4ab0c";
		wait for Clk_period;
		Addr <=  "00100001001001";
		Trees_din <= x"09004f04";
		wait for Clk_period;
		Addr <=  "00100001001010";
		Trees_din <= x"ffe32185";
		wait for Clk_period;
		Addr <=  "00100001001011";
		Trees_din <= x"11023204";
		wait for Clk_period;
		Addr <=  "00100001001100";
		Trees_din <= x"00b02185";
		wait for Clk_period;
		Addr <=  "00100001001101";
		Trees_din <= x"000a2185";
		wait for Clk_period;
		Addr <=  "00100001001110";
		Trees_din <= x"0211fd20";
		wait for Clk_period;
		Addr <=  "00100001001111";
		Trees_din <= x"08001510";
		wait for Clk_period;
		Addr <=  "00100001010000";
		Trees_din <= x"06f7d008";
		wait for Clk_period;
		Addr <=  "00100001010001";
		Trees_din <= x"0d016b04";
		wait for Clk_period;
		Addr <=  "00100001010010";
		Trees_din <= x"00102185";
		wait for Clk_period;
		Addr <=  "00100001010011";
		Trees_din <= x"ffa62185";
		wait for Clk_period;
		Addr <=  "00100001010100";
		Trees_din <= x"0afb0704";
		wait for Clk_period;
		Addr <=  "00100001010101";
		Trees_din <= x"00632185";
		wait for Clk_period;
		Addr <=  "00100001010110";
		Trees_din <= x"ffe42185";
		wait for Clk_period;
		Addr <=  "00100001010111";
		Trees_din <= x"08002608";
		wait for Clk_period;
		Addr <=  "00100001011000";
		Trees_din <= x"13fdbb04";
		wait for Clk_period;
		Addr <=  "00100001011001";
		Trees_din <= x"ffc92185";
		wait for Clk_period;
		Addr <=  "00100001011010";
		Trees_din <= x"007b2185";
		wait for Clk_period;
		Addr <=  "00100001011011";
		Trees_din <= x"0800b404";
		wait for Clk_period;
		Addr <=  "00100001011100";
		Trees_din <= x"ffeb2185";
		wait for Clk_period;
		Addr <=  "00100001011101";
		Trees_din <= x"00072185";
		wait for Clk_period;
		Addr <=  "00100001011110";
		Trees_din <= x"0af89204";
		wait for Clk_period;
		Addr <=  "00100001011111";
		Trees_din <= x"fff22185";
		wait for Clk_period;
		Addr <=  "00100001100000";
		Trees_din <= x"00742185";
		wait for Clk_period;
		Addr <=  "00100001100001";
		Trees_din <= x"02fce404";
		wait for Clk_period;
		Addr <=  "00100001100010";
		Trees_din <= x"ff9a2261";
		wait for Clk_period;
		Addr <=  "00100001100011";
		Trees_din <= x"0c02073c";
		wait for Clk_period;
		Addr <=  "00100001100100";
		Trees_din <= x"08029f20";
		wait for Clk_period;
		Addr <=  "00100001100101";
		Trees_din <= x"09005610";
		wait for Clk_period;
		Addr <=  "00100001100110";
		Trees_din <= x"0201b308";
		wait for Clk_period;
		Addr <=  "00100001100111";
		Trees_din <= x"1702f904";
		wait for Clk_period;
		Addr <=  "00100001101000";
		Trees_din <= x"ff8c2261";
		wait for Clk_period;
		Addr <=  "00100001101001";
		Trees_din <= x"00102261";
		wait for Clk_period;
		Addr <=  "00100001101010";
		Trees_din <= x"0bf96204";
		wait for Clk_period;
		Addr <=  "00100001101011";
		Trees_din <= x"00622261";
		wait for Clk_period;
		Addr <=  "00100001101100";
		Trees_din <= x"00132261";
		wait for Clk_period;
		Addr <=  "00100001101101";
		Trees_din <= x"09005608";
		wait for Clk_period;
		Addr <=  "00100001101110";
		Trees_din <= x"1d004a04";
		wait for Clk_period;
		Addr <=  "00100001101111";
		Trees_din <= x"ff492261";
		wait for Clk_period;
		Addr <=  "00100001110000";
		Trees_din <= x"ffef2261";
		wait for Clk_period;
		Addr <=  "00100001110001";
		Trees_din <= x"10048904";
		wait for Clk_period;
		Addr <=  "00100001110010";
		Trees_din <= x"000e2261";
		wait for Clk_period;
		Addr <=  "00100001110011";
		Trees_din <= x"ffb42261";
		wait for Clk_period;
		Addr <=  "00100001110100";
		Trees_din <= x"1a00e30c";
		wait for Clk_period;
		Addr <=  "00100001110101";
		Trees_din <= x"09004f04";
		wait for Clk_period;
		Addr <=  "00100001110110";
		Trees_din <= x"002e2261";
		wait for Clk_period;
		Addr <=  "00100001110111";
		Trees_din <= x"01ffc504";
		wait for Clk_period;
		Addr <=  "00100001111000";
		Trees_din <= x"00132261";
		wait for Clk_period;
		Addr <=  "00100001111001";
		Trees_din <= x"ff512261";
		wait for Clk_period;
		Addr <=  "00100001111010";
		Trees_din <= x"03fa5a08";
		wait for Clk_period;
		Addr <=  "00100001111011";
		Trees_din <= x"1f000004";
		wait for Clk_period;
		Addr <=  "00100001111100";
		Trees_din <= x"ffe62261";
		wait for Clk_period;
		Addr <=  "00100001111101";
		Trees_din <= x"ff912261";
		wait for Clk_period;
		Addr <=  "00100001111110";
		Trees_din <= x"02025304";
		wait for Clk_period;
		Addr <=  "00100001111111";
		Trees_din <= x"ffa62261";
		wait for Clk_period;
		Addr <=  "00100010000000";
		Trees_din <= x"00682261";
		wait for Clk_period;
		Addr <=  "00100010000001";
		Trees_din <= x"09004c10";
		wait for Clk_period;
		Addr <=  "00100010000010";
		Trees_din <= x"0efd5a04";
		wait for Clk_period;
		Addr <=  "00100010000011";
		Trees_din <= x"002d2261";
		wait for Clk_period;
		Addr <=  "00100010000100";
		Trees_din <= x"18004404";
		wait for Clk_period;
		Addr <=  "00100010000101";
		Trees_din <= x"ff732261";
		wait for Clk_period;
		Addr <=  "00100010000110";
		Trees_din <= x"1a00b804";
		wait for Clk_period;
		Addr <=  "00100010000111";
		Trees_din <= x"ffbd2261";
		wait for Clk_period;
		Addr <=  "00100010001000";
		Trees_din <= x"003a2261";
		wait for Clk_period;
		Addr <=  "00100010001001";
		Trees_din <= x"0c02c510";
		wait for Clk_period;
		Addr <=  "00100010001010";
		Trees_din <= x"07005808";
		wait for Clk_period;
		Addr <=  "00100010001011";
		Trees_din <= x"16001204";
		wait for Clk_period;
		Addr <=  "00100010001100";
		Trees_din <= x"008c2261";
		wait for Clk_period;
		Addr <=  "00100010001101";
		Trees_din <= x"fff12261";
		wait for Clk_period;
		Addr <=  "00100010001110";
		Trees_din <= x"02029504";
		wait for Clk_period;
		Addr <=  "00100010001111";
		Trees_din <= x"fff42261";
		wait for Clk_period;
		Addr <=  "00100010010000";
		Trees_din <= x"00802261";
		wait for Clk_period;
		Addr <=  "00100010010001";
		Trees_din <= x"0afcad08";
		wait for Clk_period;
		Addr <=  "00100010010010";
		Trees_din <= x"0208db04";
		wait for Clk_period;
		Addr <=  "00100010010011";
		Trees_din <= x"ffab2261";
		wait for Clk_period;
		Addr <=  "00100010010100";
		Trees_din <= x"002f2261";
		wait for Clk_period;
		Addr <=  "00100010010101";
		Trees_din <= x"0f00c604";
		wait for Clk_period;
		Addr <=  "00100010010110";
		Trees_din <= x"004f2261";
		wait for Clk_period;
		Addr <=  "00100010010111";
		Trees_din <= x"ffe92261";
		wait for Clk_period;
		Addr <=  "00100010011000";
		Trees_din <= x"0406be60";
		wait for Clk_period;
		Addr <=  "00100010011001";
		Trees_din <= x"04037834";
		wait for Clk_period;
		Addr <=  "00100010011010";
		Trees_din <= x"0204751c";
		wait for Clk_period;
		Addr <=  "00100010011011";
		Trees_din <= x"07005510";
		wait for Clk_period;
		Addr <=  "00100010011100";
		Trees_din <= x"1201b908";
		wait for Clk_period;
		Addr <=  "00100010011101";
		Trees_din <= x"0c039b04";
		wait for Clk_period;
		Addr <=  "00100010011110";
		Trees_din <= x"ffa8238d";
		wait for Clk_period;
		Addr <=  "00100010011111";
		Trees_din <= x"006d238d";
		wait for Clk_period;
		Addr <=  "00100010100000";
		Trees_din <= x"17004804";
		wait for Clk_period;
		Addr <=  "00100010100001";
		Trees_din <= x"ffac238d";
		wait for Clk_period;
		Addr <=  "00100010100010";
		Trees_din <= x"006d238d";
		wait for Clk_period;
		Addr <=  "00100010100011";
		Trees_din <= x"0803b608";
		wait for Clk_period;
		Addr <=  "00100010100100";
		Trees_din <= x"13f93704";
		wait for Clk_period;
		Addr <=  "00100010100101";
		Trees_din <= x"001b238d";
		wait for Clk_period;
		Addr <=  "00100010100110";
		Trees_din <= x"ff9c238d";
		wait for Clk_period;
		Addr <=  "00100010100111";
		Trees_din <= x"0070238d";
		wait for Clk_period;
		Addr <=  "00100010101000";
		Trees_din <= x"06f00008";
		wait for Clk_period;
		Addr <=  "00100010101001";
		Trees_din <= x"0009b104";
		wait for Clk_period;
		Addr <=  "00100010101010";
		Trees_din <= x"0034238d";
		wait for Clk_period;
		Addr <=  "00100010101011";
		Trees_din <= x"ff82238d";
		wait for Clk_period;
		Addr <=  "00100010101100";
		Trees_din <= x"11044408";
		wait for Clk_period;
		Addr <=  "00100010101101";
		Trees_din <= x"0e025a04";
		wait for Clk_period;
		Addr <=  "00100010101110";
		Trees_din <= x"000f238d";
		wait for Clk_period;
		Addr <=  "00100010101111";
		Trees_din <= x"ffd7238d";
		wait for Clk_period;
		Addr <=  "00100010110000";
		Trees_din <= x"11046d04";
		wait for Clk_period;
		Addr <=  "00100010110001";
		Trees_din <= x"0084238d";
		wait for Clk_period;
		Addr <=  "00100010110010";
		Trees_din <= x"ffff238d";
		wait for Clk_period;
		Addr <=  "00100010110011";
		Trees_din <= x"0b04c120";
		wait for Clk_period;
		Addr <=  "00100010110100";
		Trees_din <= x"0bfb1410";
		wait for Clk_period;
		Addr <=  "00100010110101";
		Trees_din <= x"1201de08";
		wait for Clk_period;
		Addr <=  "00100010110110";
		Trees_din <= x"1d003e04";
		wait for Clk_period;
		Addr <=  "00100010110111";
		Trees_din <= x"ffe3238d";
		wait for Clk_period;
		Addr <=  "00100010111000";
		Trees_din <= x"00bd238d";
		wait for Clk_period;
		Addr <=  "00100010111001";
		Trees_din <= x"0c01df04";
		wait for Clk_period;
		Addr <=  "00100010111010";
		Trees_din <= x"0050238d";
		wait for Clk_period;
		Addr <=  "00100010111011";
		Trees_din <= x"ff9a238d";
		wait for Clk_period;
		Addr <=  "00100010111100";
		Trees_din <= x"16023508";
		wait for Clk_period;
		Addr <=  "00100010111101";
		Trees_din <= x"1d004e04";
		wait for Clk_period;
		Addr <=  "00100010111110";
		Trees_din <= x"003a238d";
		wait for Clk_period;
		Addr <=  "00100010111111";
		Trees_din <= x"ff94238d";
		wait for Clk_period;
		Addr <=  "00100011000000";
		Trees_din <= x"0f000404";
		wait for Clk_period;
		Addr <=  "00100011000001";
		Trees_din <= x"0023238d";
		wait for Clk_period;
		Addr <=  "00100011000010";
		Trees_din <= x"ff68238d";
		wait for Clk_period;
		Addr <=  "00100011000011";
		Trees_din <= x"05fdf608";
		wait for Clk_period;
		Addr <=  "00100011000100";
		Trees_din <= x"03041704";
		wait for Clk_period;
		Addr <=  "00100011000101";
		Trees_din <= x"00a5238d";
		wait for Clk_period;
		Addr <=  "00100011000110";
		Trees_din <= x"ffec238d";
		wait for Clk_period;
		Addr <=  "00100011000111";
		Trees_din <= x"ffb9238d";
		wait for Clk_period;
		Addr <=  "00100011001000";
		Trees_din <= x"1d004114";
		wait for Clk_period;
		Addr <=  "00100011001001";
		Trees_din <= x"0105650c";
		wait for Clk_period;
		Addr <=  "00100011001010";
		Trees_din <= x"02032e04";
		wait for Clk_period;
		Addr <=  "00100011001011";
		Trees_din <= x"ff95238d";
		wait for Clk_period;
		Addr <=  "00100011001100";
		Trees_din <= x"13fdca04";
		wait for Clk_period;
		Addr <=  "00100011001101";
		Trees_din <= x"0066238d";
		wait for Clk_period;
		Addr <=  "00100011001110";
		Trees_din <= x"0006238d";
		wait for Clk_period;
		Addr <=  "00100011001111";
		Trees_din <= x"14008c04";
		wait for Clk_period;
		Addr <=  "00100011010000";
		Trees_din <= x"fffb238d";
		wait for Clk_period;
		Addr <=  "00100011010001";
		Trees_din <= x"ff60238d";
		wait for Clk_period;
		Addr <=  "00100011010010";
		Trees_din <= x"1c00350c";
		wait for Clk_period;
		Addr <=  "00100011010011";
		Trees_din <= x"0b046408";
		wait for Clk_period;
		Addr <=  "00100011010100";
		Trees_din <= x"05fa9204";
		wait for Clk_period;
		Addr <=  "00100011010101";
		Trees_din <= x"00b2238d";
		wait for Clk_period;
		Addr <=  "00100011010110";
		Trees_din <= x"001b238d";
		wait for Clk_period;
		Addr <=  "00100011010111";
		Trees_din <= x"ffba238d";
		wait for Clk_period;
		Addr <=  "00100011011000";
		Trees_din <= x"0900580c";
		wait for Clk_period;
		Addr <=  "00100011011001";
		Trees_din <= x"10053b08";
		wait for Clk_period;
		Addr <=  "00100011011010";
		Trees_din <= x"040d1104";
		wait for Clk_period;
		Addr <=  "00100011011011";
		Trees_din <= x"ff84238d";
		wait for Clk_period;
		Addr <=  "00100011011100";
		Trees_din <= x"fffb238d";
		wait for Clk_period;
		Addr <=  "00100011011101";
		Trees_din <= x"002c238d";
		wait for Clk_period;
		Addr <=  "00100011011110";
		Trees_din <= x"11028408";
		wait for Clk_period;
		Addr <=  "00100011011111";
		Trees_din <= x"0202d904";
		wait for Clk_period;
		Addr <=  "00100011100000";
		Trees_din <= x"ff9b238d";
		wait for Clk_period;
		Addr <=  "00100011100001";
		Trees_din <= x"003b238d";
		wait for Clk_period;
		Addr <=  "00100011100010";
		Trees_din <= x"0064238d";
		wait for Clk_period;
		Addr <=  "00100011100011";
		Trees_din <= x"020baf74";
		wait for Clk_period;
		Addr <=  "00100011100100";
		Trees_din <= x"04f95838";
		wait for Clk_period;
		Addr <=  "00100011100101";
		Trees_din <= x"0d02541c";
		wait for Clk_period;
		Addr <=  "00100011100110";
		Trees_din <= x"0effcc10";
		wait for Clk_period;
		Addr <=  "00100011100111";
		Trees_din <= x"0a028808";
		wait for Clk_period;
		Addr <=  "00100011101000";
		Trees_din <= x"04f60a04";
		wait for Clk_period;
		Addr <=  "00100011101001";
		Trees_din <= x"000b24e1";
		wait for Clk_period;
		Addr <=  "00100011101010";
		Trees_din <= x"ff8f24e1";
		wait for Clk_period;
		Addr <=  "00100011101011";
		Trees_din <= x"04f81504";
		wait for Clk_period;
		Addr <=  "00100011101100";
		Trees_din <= x"ffe624e1";
		wait for Clk_period;
		Addr <=  "00100011101101";
		Trees_din <= x"00a824e1";
		wait for Clk_period;
		Addr <=  "00100011101110";
		Trees_din <= x"08034d08";
		wait for Clk_period;
		Addr <=  "00100011101111";
		Trees_din <= x"14002604";
		wait for Clk_period;
		Addr <=  "00100011110000";
		Trees_din <= x"000424e1";
		wait for Clk_period;
		Addr <=  "00100011110001";
		Trees_din <= x"ff6c24e1";
		wait for Clk_period;
		Addr <=  "00100011110010";
		Trees_din <= x"002b24e1";
		wait for Clk_period;
		Addr <=  "00100011110011";
		Trees_din <= x"1b003610";
		wait for Clk_period;
		Addr <=  "00100011110100";
		Trees_din <= x"0c01cf08";
		wait for Clk_period;
		Addr <=  "00100011110101";
		Trees_din <= x"13fdbe04";
		wait for Clk_period;
		Addr <=  "00100011110110";
		Trees_din <= x"00db24e1";
		wait for Clk_period;
		Addr <=  "00100011110111";
		Trees_din <= x"002024e1";
		wait for Clk_period;
		Addr <=  "00100011111000";
		Trees_din <= x"1102c604";
		wait for Clk_period;
		Addr <=  "00100011111001";
		Trees_din <= x"ff9c24e1";
		wait for Clk_period;
		Addr <=  "00100011111010";
		Trees_din <= x"005124e1";
		wait for Clk_period;
		Addr <=  "00100011111011";
		Trees_din <= x"16001604";
		wait for Clk_period;
		Addr <=  "00100011111100";
		Trees_din <= x"006324e1";
		wait for Clk_period;
		Addr <=  "00100011111101";
		Trees_din <= x"0c016804";
		wait for Clk_period;
		Addr <=  "00100011111110";
		Trees_din <= x"001c24e1";
		wait for Clk_period;
		Addr <=  "00100011111111";
		Trees_din <= x"ff8624e1";
		wait for Clk_period;
		Addr <=  "00100100000000";
		Trees_din <= x"04fba420";
		wait for Clk_period;
		Addr <=  "00100100000001";
		Trees_din <= x"07005910";
		wait for Clk_period;
		Addr <=  "00100100000010";
		Trees_din <= x"03fee208";
		wait for Clk_period;
		Addr <=  "00100100000011";
		Trees_din <= x"06f51c04";
		wait for Clk_period;
		Addr <=  "00100100000100";
		Trees_din <= x"003824e1";
		wait for Clk_period;
		Addr <=  "00100100000101";
		Trees_din <= x"ffbe24e1";
		wait for Clk_period;
		Addr <=  "00100100000110";
		Trees_din <= x"02024904";
		wait for Clk_period;
		Addr <=  "00100100000111";
		Trees_din <= x"ffd224e1";
		wait for Clk_period;
		Addr <=  "00100100001000";
		Trees_din <= x"008224e1";
		wait for Clk_period;
		Addr <=  "00100100001001";
		Trees_din <= x"10028508";
		wait for Clk_period;
		Addr <=  "00100100001010";
		Trees_din <= x"000f3604";
		wait for Clk_period;
		Addr <=  "00100100001011";
		Trees_din <= x"000724e1";
		wait for Clk_period;
		Addr <=  "00100100001100";
		Trees_din <= x"ffa124e1";
		wait for Clk_period;
		Addr <=  "00100100001101";
		Trees_din <= x"02039104";
		wait for Clk_period;
		Addr <=  "00100100001110";
		Trees_din <= x"001424e1";
		wait for Clk_period;
		Addr <=  "00100100001111";
		Trees_din <= x"00c024e1";
		wait for Clk_period;
		Addr <=  "00100100010000";
		Trees_din <= x"0c00460c";
		wait for Clk_period;
		Addr <=  "00100100010001";
		Trees_din <= x"1d004004";
		wait for Clk_period;
		Addr <=  "00100100010010";
		Trees_din <= x"003724e1";
		wait for Clk_period;
		Addr <=  "00100100010011";
		Trees_din <= x"01fc0b04";
		wait for Clk_period;
		Addr <=  "00100100010100";
		Trees_din <= x"002824e1";
		wait for Clk_period;
		Addr <=  "00100100010101";
		Trees_din <= x"ff7724e1";
		wait for Clk_period;
		Addr <=  "00100100010110";
		Trees_din <= x"1603f908";
		wait for Clk_period;
		Addr <=  "00100100010111";
		Trees_din <= x"0e02f104";
		wait for Clk_period;
		Addr <=  "00100100011000";
		Trees_din <= x"fff124e1";
		wait for Clk_period;
		Addr <=  "00100100011001";
		Trees_din <= x"002824e1";
		wait for Clk_period;
		Addr <=  "00100100011010";
		Trees_din <= x"1a00db04";
		wait for Clk_period;
		Addr <=  "00100100011011";
		Trees_din <= x"007b24e1";
		wait for Clk_period;
		Addr <=  "00100100011100";
		Trees_din <= x"ffd824e1";
		wait for Clk_period;
		Addr <=  "00100100011101";
		Trees_din <= x"0001c404";
		wait for Clk_period;
		Addr <=  "00100100011110";
		Trees_din <= x"007e24e1";
		wait for Clk_period;
		Addr <=  "00100100011111";
		Trees_din <= x"06f34c18";
		wait for Clk_period;
		Addr <=  "00100100100000";
		Trees_din <= x"01025908";
		wait for Clk_period;
		Addr <=  "00100100100001";
		Trees_din <= x"0afc3704";
		wait for Clk_period;
		Addr <=  "00100100100010";
		Trees_din <= x"ff3524e1";
		wait for Clk_period;
		Addr <=  "00100100100011";
		Trees_din <= x"fff024e1";
		wait for Clk_period;
		Addr <=  "00100100100100";
		Trees_din <= x"05fc5d08";
		wait for Clk_period;
		Addr <=  "00100100100101";
		Trees_din <= x"1201da04";
		wait for Clk_period;
		Addr <=  "00100100100110";
		Trees_din <= x"001c24e1";
		wait for Clk_period;
		Addr <=  "00100100100111";
		Trees_din <= x"ffa924e1";
		wait for Clk_period;
		Addr <=  "00100100101000";
		Trees_din <= x"0c01ad04";
		wait for Clk_period;
		Addr <=  "00100100101001";
		Trees_din <= x"007d24e1";
		wait for Clk_period;
		Addr <=  "00100100101010";
		Trees_din <= x"000c24e1";
		wait for Clk_period;
		Addr <=  "00100100101011";
		Trees_din <= x"07005a0c";
		wait for Clk_period;
		Addr <=  "00100100101100";
		Trees_din <= x"08035608";
		wait for Clk_period;
		Addr <=  "00100100101101";
		Trees_din <= x"14031e04";
		wait for Clk_period;
		Addr <=  "00100100101110";
		Trees_din <= x"005c24e1";
		wait for Clk_period;
		Addr <=  "00100100101111";
		Trees_din <= x"ffff24e1";
		wait for Clk_period;
		Addr <=  "00100100110000";
		Trees_din <= x"ffaf24e1";
		wait for Clk_period;
		Addr <=  "00100100110001";
		Trees_din <= x"0afb1508";
		wait for Clk_period;
		Addr <=  "00100100110010";
		Trees_din <= x"0b03e304";
		wait for Clk_period;
		Addr <=  "00100100110011";
		Trees_din <= x"ff7424e1";
		wait for Clk_period;
		Addr <=  "00100100110100";
		Trees_din <= x"000724e1";
		wait for Clk_period;
		Addr <=  "00100100110101";
		Trees_din <= x"19008b04";
		wait for Clk_period;
		Addr <=  "00100100110110";
		Trees_din <= x"001424e1";
		wait for Clk_period;
		Addr <=  "00100100110111";
		Trees_din <= x"005224e1";
		wait for Clk_period;
		Addr <=  "00100100111000";
		Trees_din <= x"0c020760";
		wait for Clk_period;
		Addr <=  "00100100111001";
		Trees_din <= x"08029f38";
		wait for Clk_period;
		Addr <=  "00100100111010";
		Trees_din <= x"0406be20";
		wait for Clk_period;
		Addr <=  "00100100111011";
		Trees_din <= x"1c002f10";
		wait for Clk_period;
		Addr <=  "00100100111100";
		Trees_din <= x"0201e308";
		wait for Clk_period;
		Addr <=  "00100100111101";
		Trees_din <= x"04032b04";
		wait for Clk_period;
		Addr <=  "00100100111110";
		Trees_din <= x"ff8a2635";
		wait for Clk_period;
		Addr <=  "00100100111111";
		Trees_din <= x"00262635";
		wait for Clk_period;
		Addr <=  "00100101000000";
		Trees_din <= x"05f9ab04";
		wait for Clk_period;
		Addr <=  "00100101000001";
		Trees_din <= x"ffe72635";
		wait for Clk_period;
		Addr <=  "00100101000010";
		Trees_din <= x"004b2635";
		wait for Clk_period;
		Addr <=  "00100101000011";
		Trees_din <= x"1c003108";
		wait for Clk_period;
		Addr <=  "00100101000100";
		Trees_din <= x"13004104";
		wait for Clk_period;
		Addr <=  "00100101000101";
		Trees_din <= x"ff7e2635";
		wait for Clk_period;
		Addr <=  "00100101000110";
		Trees_din <= x"00352635";
		wait for Clk_period;
		Addr <=  "00100101000111";
		Trees_din <= x"03fa4604";
		wait for Clk_period;
		Addr <=  "00100101001000";
		Trees_din <= x"ffdd2635";
		wait for Clk_period;
		Addr <=  "00100101001001";
		Trees_din <= x"001e2635";
		wait for Clk_period;
		Addr <=  "00100101001010";
		Trees_din <= x"00fd640c";
		wait for Clk_period;
		Addr <=  "00100101001011";
		Trees_din <= x"0202d904";
		wait for Clk_period;
		Addr <=  "00100101001100";
		Trees_din <= x"ffb32635";
		wait for Clk_period;
		Addr <=  "00100101001101";
		Trees_din <= x"05fa9204";
		wait for Clk_period;
		Addr <=  "00100101001110";
		Trees_din <= x"00632635";
		wait for Clk_period;
		Addr <=  "00100101001111";
		Trees_din <= x"ffd12635";
		wait for Clk_period;
		Addr <=  "00100101010000";
		Trees_din <= x"1703c808";
		wait for Clk_period;
		Addr <=  "00100101010001";
		Trees_din <= x"01ffe604";
		wait for Clk_period;
		Addr <=  "00100101010010";
		Trees_din <= x"ffe42635";
		wait for Clk_period;
		Addr <=  "00100101010011";
		Trees_din <= x"ff672635";
		wait for Clk_period;
		Addr <=  "00100101010100";
		Trees_din <= x"00252635";
		wait for Clk_period;
		Addr <=  "00100101010101";
		Trees_din <= x"03fe2518";
		wait for Clk_period;
		Addr <=  "00100101010110";
		Trees_din <= x"0700540c";
		wait for Clk_period;
		Addr <=  "00100101010111";
		Trees_din <= x"02083204";
		wait for Clk_period;
		Addr <=  "00100101011000";
		Trees_din <= x"ff8a2635";
		wait for Clk_period;
		Addr <=  "00100101011001";
		Trees_din <= x"07005004";
		wait for Clk_period;
		Addr <=  "00100101011010";
		Trees_din <= x"00132635";
		wait for Clk_period;
		Addr <=  "00100101011011";
		Trees_din <= x"005a2635";
		wait for Clk_period;
		Addr <=  "00100101011100";
		Trees_din <= x"05f9bd04";
		wait for Clk_period;
		Addr <=  "00100101011101";
		Trees_din <= x"ffe52635";
		wait for Clk_period;
		Addr <=  "00100101011110";
		Trees_din <= x"0d008304";
		wait for Clk_period;
		Addr <=  "00100101011111";
		Trees_din <= x"ffd52635";
		wait for Clk_period;
		Addr <=  "00100101100000";
		Trees_din <= x"ff592635";
		wait for Clk_period;
		Addr <=  "00100101100001";
		Trees_din <= x"15009e08";
		wait for Clk_period;
		Addr <=  "00100101100010";
		Trees_din <= x"0101d104";
		wait for Clk_period;
		Addr <=  "00100101100011";
		Trees_din <= x"00092635";
		wait for Clk_period;
		Addr <=  "00100101100100";
		Trees_din <= x"ffa42635";
		wait for Clk_period;
		Addr <=  "00100101100101";
		Trees_din <= x"06f50b04";
		wait for Clk_period;
		Addr <=  "00100101100110";
		Trees_din <= x"006a2635";
		wait for Clk_period;
		Addr <=  "00100101100111";
		Trees_din <= x"fffb2635";
		wait for Clk_period;
		Addr <=  "00100101101000";
		Trees_din <= x"09004c10";
		wait for Clk_period;
		Addr <=  "00100101101001";
		Trees_din <= x"12028508";
		wait for Clk_period;
		Addr <=  "00100101101010";
		Trees_din <= x"0d037304";
		wait for Clk_period;
		Addr <=  "00100101101011";
		Trees_din <= x"ff7a2635";
		wait for Clk_period;
		Addr <=  "00100101101100";
		Trees_din <= x"ffdb2635";
		wait for Clk_period;
		Addr <=  "00100101101101";
		Trees_din <= x"17001c04";
		wait for Clk_period;
		Addr <=  "00100101101110";
		Trees_din <= x"ffb92635";
		wait for Clk_period;
		Addr <=  "00100101101111";
		Trees_din <= x"00452635";
		wait for Clk_period;
		Addr <=  "00100101110000";
		Trees_din <= x"0c02c51c";
		wait for Clk_period;
		Addr <=  "00100101110001";
		Trees_din <= x"07005910";
		wait for Clk_period;
		Addr <=  "00100101110010";
		Trees_din <= x"16006908";
		wait for Clk_period;
		Addr <=  "00100101110011";
		Trees_din <= x"0206a304";
		wait for Clk_period;
		Addr <=  "00100101110100";
		Trees_din <= x"00992635";
		wait for Clk_period;
		Addr <=  "00100101110101";
		Trees_din <= x"ffed2635";
		wait for Clk_period;
		Addr <=  "00100101110110";
		Trees_din <= x"0209bd04";
		wait for Clk_period;
		Addr <=  "00100101110111";
		Trees_din <= x"ffdc2635";
		wait for Clk_period;
		Addr <=  "00100101111000";
		Trees_din <= x"00552635";
		wait for Clk_period;
		Addr <=  "00100101111001";
		Trees_din <= x"0202ac04";
		wait for Clk_period;
		Addr <=  "00100101111010";
		Trees_din <= x"ffed2635";
		wait for Clk_period;
		Addr <=  "00100101111011";
		Trees_din <= x"0f032a04";
		wait for Clk_period;
		Addr <=  "00100101111100";
		Trees_din <= x"008d2635";
		wait for Clk_period;
		Addr <=  "00100101111101";
		Trees_din <= x"000c2635";
		wait for Clk_period;
		Addr <=  "00100101111110";
		Trees_din <= x"04001f10";
		wait for Clk_period;
		Addr <=  "00100101111111";
		Trees_din <= x"02085c08";
		wait for Clk_period;
		Addr <=  "00100110000000";
		Trees_din <= x"06f87f04";
		wait for Clk_period;
		Addr <=  "00100110000001";
		Trees_din <= x"ff972635";
		wait for Clk_period;
		Addr <=  "00100110000010";
		Trees_din <= x"000e2635";
		wait for Clk_period;
		Addr <=  "00100110000011";
		Trees_din <= x"04fea404";
		wait for Clk_period;
		Addr <=  "00100110000100";
		Trees_din <= x"00382635";
		wait for Clk_period;
		Addr <=  "00100110000101";
		Trees_din <= x"ff942635";
		wait for Clk_period;
		Addr <=  "00100110000110";
		Trees_din <= x"12013b08";
		wait for Clk_period;
		Addr <=  "00100110000111";
		Trees_din <= x"13fdda04";
		wait for Clk_period;
		Addr <=  "00100110001000";
		Trees_din <= x"00122635";
		wait for Clk_period;
		Addr <=  "00100110001001";
		Trees_din <= x"00862635";
		wait for Clk_period;
		Addr <=  "00100110001010";
		Trees_din <= x"03fd6504";
		wait for Clk_period;
		Addr <=  "00100110001011";
		Trees_din <= x"00252635";
		wait for Clk_period;
		Addr <=  "00100110001100";
		Trees_din <= x"ffb22635";
		wait for Clk_period;
		Addr <=  "00100110001101";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00100110001110";
		Trees_din <= x"0211fd60";
		wait for Clk_period;
		Addr <=  "00100110001111";
		Trees_din <= x"1b002e24";
		wait for Clk_period;
		Addr <=  "00100110010000";
		Trees_din <= x"21000018";
		wait for Clk_period;
		Addr <=  "00100110010001";
		Trees_din <= x"1d003c10";
		wait for Clk_period;
		Addr <=  "00100110010010";
		Trees_din <= x"1d003608";
		wait for Clk_period;
		Addr <=  "00100110010011";
		Trees_din <= x"13fe6b04";
		wait for Clk_period;
		Addr <=  "00100110010100";
		Trees_din <= x"003a2705";
		wait for Clk_period;
		Addr <=  "00100110010101";
		Trees_din <= x"ffbf2705";
		wait for Clk_period;
		Addr <=  "00100110010110";
		Trees_din <= x"12000f04";
		wait for Clk_period;
		Addr <=  "00100110010111";
		Trees_din <= x"fff12705";
		wait for Clk_period;
		Addr <=  "00100110011000";
		Trees_din <= x"ff882705";
		wait for Clk_period;
		Addr <=  "00100110011001";
		Trees_din <= x"09005004";
		wait for Clk_period;
		Addr <=  "00100110011010";
		Trees_din <= x"005d2705";
		wait for Clk_period;
		Addr <=  "00100110011011";
		Trees_din <= x"00112705";
		wait for Clk_period;
		Addr <=  "00100110011100";
		Trees_din <= x"1900a704";
		wait for Clk_period;
		Addr <=  "00100110011101";
		Trees_din <= x"ffc22705";
		wait for Clk_period;
		Addr <=  "00100110011110";
		Trees_din <= x"18003604";
		wait for Clk_period;
		Addr <=  "00100110011111";
		Trees_din <= x"007e2705";
		wait for Clk_period;
		Addr <=  "00100110100000";
		Trees_din <= x"00042705";
		wait for Clk_period;
		Addr <=  "00100110100001";
		Trees_din <= x"1e006020";
		wait for Clk_period;
		Addr <=  "00100110100010";
		Trees_din <= x"1d003f10";
		wait for Clk_period;
		Addr <=  "00100110100011";
		Trees_din <= x"12011f08";
		wait for Clk_period;
		Addr <=  "00100110100100";
		Trees_din <= x"0f000404";
		wait for Clk_period;
		Addr <=  "00100110100101";
		Trees_din <= x"00592705";
		wait for Clk_period;
		Addr <=  "00100110100110";
		Trees_din <= x"ffbc2705";
		wait for Clk_period;
		Addr <=  "00100110100111";
		Trees_din <= x"04025d04";
		wait for Clk_period;
		Addr <=  "00100110101000";
		Trees_din <= x"004d2705";
		wait for Clk_period;
		Addr <=  "00100110101001";
		Trees_din <= x"ffd72705";
		wait for Clk_period;
		Addr <=  "00100110101010";
		Trees_din <= x"0c022408";
		wait for Clk_period;
		Addr <=  "00100110101011";
		Trees_din <= x"0eff8004";
		wait for Clk_period;
		Addr <=  "00100110101100";
		Trees_din <= x"ff9f2705";
		wait for Clk_period;
		Addr <=  "00100110101101";
		Trees_din <= x"005c2705";
		wait for Clk_period;
		Addr <=  "00100110101110";
		Trees_din <= x"0a01b504";
		wait for Clk_period;
		Addr <=  "00100110101111";
		Trees_din <= x"002c2705";
		wait for Clk_period;
		Addr <=  "00100110110000";
		Trees_din <= x"00ae2705";
		wait for Clk_period;
		Addr <=  "00100110110001";
		Trees_din <= x"1e00620c";
		wait for Clk_period;
		Addr <=  "00100110110010";
		Trees_din <= x"1500a708";
		wait for Clk_period;
		Addr <=  "00100110110011";
		Trees_din <= x"17000204";
		wait for Clk_period;
		Addr <=  "00100110110100";
		Trees_din <= x"ffec2705";
		wait for Clk_period;
		Addr <=  "00100110110101";
		Trees_din <= x"ff5c2705";
		wait for Clk_period;
		Addr <=  "00100110110110";
		Trees_din <= x"00462705";
		wait for Clk_period;
		Addr <=  "00100110110111";
		Trees_din <= x"0800b708";
		wait for Clk_period;
		Addr <=  "00100110111000";
		Trees_din <= x"0a016304";
		wait for Clk_period;
		Addr <=  "00100110111001";
		Trees_din <= x"00022705";
		wait for Clk_period;
		Addr <=  "00100110111010";
		Trees_din <= x"ffbd2705";
		wait for Clk_period;
		Addr <=  "00100110111011";
		Trees_din <= x"06fb2904";
		wait for Clk_period;
		Addr <=  "00100110111100";
		Trees_din <= x"00162705";
		wait for Clk_period;
		Addr <=  "00100110111101";
		Trees_din <= x"ffa42705";
		wait for Clk_period;
		Addr <=  "00100110111110";
		Trees_din <= x"17034f04";
		wait for Clk_period;
		Addr <=  "00100110111111";
		Trees_din <= x"00642705";
		wait for Clk_period;
		Addr <=  "00100111000000";
		Trees_din <= x"ffdf2705";
		wait for Clk_period;
		Addr <=  "00100111000001";
		Trees_din <= x"0207142c";
		wait for Clk_period;
		Addr <=  "00100111000010";
		Trees_din <= x"0c003208";
		wait for Clk_period;
		Addr <=  "00100111000011";
		Trees_din <= x"06f96104";
		wait for Clk_period;
		Addr <=  "00100111000100";
		Trees_din <= x"ff872799";
		wait for Clk_period;
		Addr <=  "00100111000101";
		Trees_din <= x"00182799";
		wait for Clk_period;
		Addr <=  "00100111000110";
		Trees_din <= x"0af7a504";
		wait for Clk_period;
		Addr <=  "00100111000111";
		Trees_din <= x"ff9b2799";
		wait for Clk_period;
		Addr <=  "00100111001000";
		Trees_din <= x"1702f910";
		wait for Clk_period;
		Addr <=  "00100111001001";
		Trees_din <= x"1603b408";
		wait for Clk_period;
		Addr <=  "00100111001010";
		Trees_din <= x"1d003e04";
		wait for Clk_period;
		Addr <=  "00100111001011";
		Trees_din <= x"ffd82799";
		wait for Clk_period;
		Addr <=  "00100111001100";
		Trees_din <= x"00112799";
		wait for Clk_period;
		Addr <=  "00100111001101";
		Trees_din <= x"1500ac04";
		wait for Clk_period;
		Addr <=  "00100111001110";
		Trees_din <= x"ff932799";
		wait for Clk_period;
		Addr <=  "00100111001111";
		Trees_din <= x"00412799";
		wait for Clk_period;
		Addr <=  "00100111010000";
		Trees_din <= x"0f000c08";
		wait for Clk_period;
		Addr <=  "00100111010001";
		Trees_din <= x"13f90804";
		wait for Clk_period;
		Addr <=  "00100111010010";
		Trees_din <= x"00142799";
		wait for Clk_period;
		Addr <=  "00100111010011";
		Trees_din <= x"00892799";
		wait for Clk_period;
		Addr <=  "00100111010100";
		Trees_din <= x"04007b04";
		wait for Clk_period;
		Addr <=  "00100111010101";
		Trees_din <= x"ffac2799";
		wait for Clk_period;
		Addr <=  "00100111010110";
		Trees_din <= x"003a2799";
		wait for Clk_period;
		Addr <=  "00100111010111";
		Trees_din <= x"08000108";
		wait for Clk_period;
		Addr <=  "00100111011000";
		Trees_din <= x"15008004";
		wait for Clk_period;
		Addr <=  "00100111011001";
		Trees_din <= x"00042799";
		wait for Clk_period;
		Addr <=  "00100111011010";
		Trees_din <= x"007e2799";
		wait for Clk_period;
		Addr <=  "00100111011011";
		Trees_din <= x"10068314";
		wait for Clk_period;
		Addr <=  "00100111011100";
		Trees_din <= x"03048810";
		wait for Clk_period;
		Addr <=  "00100111011101";
		Trees_din <= x"10057f08";
		wait for Clk_period;
		Addr <=  "00100111011110";
		Trees_din <= x"02077504";
		wait for Clk_period;
		Addr <=  "00100111011111";
		Trees_din <= x"00472799";
		wait for Clk_period;
		Addr <=  "00100111100000";
		Trees_din <= x"ffff2799";
		wait for Clk_period;
		Addr <=  "00100111100001";
		Trees_din <= x"04ffda04";
		wait for Clk_period;
		Addr <=  "00100111100010";
		Trees_din <= x"ffb12799";
		wait for Clk_period;
		Addr <=  "00100111100011";
		Trees_din <= x"00542799";
		wait for Clk_period;
		Addr <=  "00100111100100";
		Trees_din <= x"00712799";
		wait for Clk_period;
		Addr <=  "00100111100101";
		Trees_din <= x"00742799";
		wait for Clk_period;
		Addr <=  "00100111100110";
		Trees_din <= x"02083250";
		wait for Clk_period;
		Addr <=  "00100111100111";
		Trees_din <= x"1b00452c";
		wait for Clk_period;
		Addr <=  "00100111101000";
		Trees_din <= x"18004618";
		wait for Clk_period;
		Addr <=  "00100111101001";
		Trees_din <= x"1d00470c";
		wait for Clk_period;
		Addr <=  "00100111101010";
		Trees_din <= x"01107308";
		wait for Clk_period;
		Addr <=  "00100111101011";
		Trees_din <= x"1d003d04";
		wait for Clk_period;
		Addr <=  "00100111101100";
		Trees_din <= x"ffe928a5";
		wait for Clk_period;
		Addr <=  "00100111101101";
		Trees_din <= x"001e28a5";
		wait for Clk_period;
		Addr <=  "00100111101110";
		Trees_din <= x"ff8928a5";
		wait for Clk_period;
		Addr <=  "00100111101111";
		Trees_din <= x"15008f04";
		wait for Clk_period;
		Addr <=  "00100111110000";
		Trees_din <= x"005028a5";
		wait for Clk_period;
		Addr <=  "00100111110001";
		Trees_din <= x"0e039c04";
		wait for Clk_period;
		Addr <=  "00100111110010";
		Trees_din <= x"ff7128a5";
		wait for Clk_period;
		Addr <=  "00100111110011";
		Trees_din <= x"000a28a5";
		wait for Clk_period;
		Addr <=  "00100111110100";
		Trees_din <= x"10f77408";
		wait for Clk_period;
		Addr <=  "00100111110101";
		Trees_din <= x"0204f604";
		wait for Clk_period;
		Addr <=  "00100111110110";
		Trees_din <= x"ffe828a5";
		wait for Clk_period;
		Addr <=  "00100111110111";
		Trees_din <= x"00a728a5";
		wait for Clk_period;
		Addr <=  "00100111111000";
		Trees_din <= x"0f000204";
		wait for Clk_period;
		Addr <=  "00100111111001";
		Trees_din <= x"003b28a5";
		wait for Clk_period;
		Addr <=  "00100111111010";
		Trees_din <= x"08002d04";
		wait for Clk_period;
		Addr <=  "00100111111011";
		Trees_din <= x"000e28a5";
		wait for Clk_period;
		Addr <=  "00100111111100";
		Trees_din <= x"ff8228a5";
		wait for Clk_period;
		Addr <=  "00100111111101";
		Trees_din <= x"06f84b1c";
		wait for Clk_period;
		Addr <=  "00100111111110";
		Trees_din <= x"0800ad10";
		wait for Clk_period;
		Addr <=  "00100111111111";
		Trees_din <= x"19007f08";
		wait for Clk_period;
		Addr <=  "00101000000000";
		Trees_din <= x"05fd2704";
		wait for Clk_period;
		Addr <=  "00101000000001";
		Trees_din <= x"ff8c28a5";
		wait for Clk_period;
		Addr <=  "00101000000010";
		Trees_din <= x"002c28a5";
		wait for Clk_period;
		Addr <=  "00101000000011";
		Trees_din <= x"13fdc104";
		wait for Clk_period;
		Addr <=  "00101000000100";
		Trees_din <= x"ffe028a5";
		wait for Clk_period;
		Addr <=  "00101000000101";
		Trees_din <= x"006f28a5";
		wait for Clk_period;
		Addr <=  "00101000000110";
		Trees_din <= x"10fb2504";
		wait for Clk_period;
		Addr <=  "00101000000111";
		Trees_din <= x"ffe728a5";
		wait for Clk_period;
		Addr <=  "00101000001000";
		Trees_din <= x"02039104";
		wait for Clk_period;
		Addr <=  "00101000001001";
		Trees_din <= x"001c28a5";
		wait for Clk_period;
		Addr <=  "00101000001010";
		Trees_din <= x"00ab28a5";
		wait for Clk_period;
		Addr <=  "00101000001011";
		Trees_din <= x"03011204";
		wait for Clk_period;
		Addr <=  "00101000001100";
		Trees_din <= x"ff8c28a5";
		wait for Clk_period;
		Addr <=  "00101000001101";
		Trees_din <= x"fffd28a5";
		wait for Clk_period;
		Addr <=  "00101000001110";
		Trees_din <= x"08000108";
		wait for Clk_period;
		Addr <=  "00101000001111";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00101000010000";
		Trees_din <= x"001728a5";
		wait for Clk_period;
		Addr <=  "00101000010001";
		Trees_din <= x"007e28a5";
		wait for Clk_period;
		Addr <=  "00101000010010";
		Trees_din <= x"000d6314";
		wait for Clk_period;
		Addr <=  "00101000010011";
		Trees_din <= x"04f69f04";
		wait for Clk_period;
		Addr <=  "00101000010100";
		Trees_din <= x"007a28a5";
		wait for Clk_period;
		Addr <=  "00101000010101";
		Trees_din <= x"0a03e208";
		wait for Clk_period;
		Addr <=  "00101000010110";
		Trees_din <= x"06f98d04";
		wait for Clk_period;
		Addr <=  "00101000010111";
		Trees_din <= x"002128a5";
		wait for Clk_period;
		Addr <=  "00101000011000";
		Trees_din <= x"ffbb28a5";
		wait for Clk_period;
		Addr <=  "00101000011001";
		Trees_din <= x"0bf9f604";
		wait for Clk_period;
		Addr <=  "00101000011010";
		Trees_din <= x"ff7228a5";
		wait for Clk_period;
		Addr <=  "00101000011011";
		Trees_din <= x"001d28a5";
		wait for Clk_period;
		Addr <=  "00101000011100";
		Trees_din <= x"08022010";
		wait for Clk_period;
		Addr <=  "00101000011101";
		Trees_din <= x"0f00ba08";
		wait for Clk_period;
		Addr <=  "00101000011110";
		Trees_din <= x"16037104";
		wait for Clk_period;
		Addr <=  "00101000011111";
		Trees_din <= x"004228a5";
		wait for Clk_period;
		Addr <=  "00101000100000";
		Trees_din <= x"ffd328a5";
		wait for Clk_period;
		Addr <=  "00101000100001";
		Trees_din <= x"1c002904";
		wait for Clk_period;
		Addr <=  "00101000100010";
		Trees_din <= x"001928a5";
		wait for Clk_period;
		Addr <=  "00101000100011";
		Trees_din <= x"ff9928a5";
		wait for Clk_period;
		Addr <=  "00101000100100";
		Trees_din <= x"09005004";
		wait for Clk_period;
		Addr <=  "00101000100101";
		Trees_din <= x"ffcb28a5";
		wait for Clk_period;
		Addr <=  "00101000100110";
		Trees_din <= x"12027604";
		wait for Clk_period;
		Addr <=  "00101000100111";
		Trees_din <= x"008228a5";
		wait for Clk_period;
		Addr <=  "00101000101000";
		Trees_din <= x"000828a5";
		wait for Clk_period;
		Addr <=  "00101000101001";
		Trees_din <= x"1104aa54";
		wait for Clk_period;
		Addr <=  "00101000101010";
		Trees_din <= x"1103b928";
		wait for Clk_period;
		Addr <=  "00101000101011";
		Trees_din <= x"07005e20";
		wait for Clk_period;
		Addr <=  "00101000101100";
		Trees_din <= x"0c006e10";
		wait for Clk_period;
		Addr <=  "00101000101101";
		Trees_din <= x"0c006108";
		wait for Clk_period;
		Addr <=  "00101000101110";
		Trees_din <= x"10027704";
		wait for Clk_period;
		Addr <=  "00101000101111";
		Trees_din <= x"ff9f2961";
		wait for Clk_period;
		Addr <=  "00101000110000";
		Trees_din <= x"00212961";
		wait for Clk_period;
		Addr <=  "00101000110001";
		Trees_din <= x"15009b04";
		wait for Clk_period;
		Addr <=  "00101000110010";
		Trees_din <= x"00842961";
		wait for Clk_period;
		Addr <=  "00101000110011";
		Trees_din <= x"00112961";
		wait for Clk_period;
		Addr <=  "00101000110100";
		Trees_din <= x"0c00ad08";
		wait for Clk_period;
		Addr <=  "00101000110101";
		Trees_din <= x"06f4d304";
		wait for Clk_period;
		Addr <=  "00101000110110";
		Trees_din <= x"ff7c2961";
		wait for Clk_period;
		Addr <=  "00101000110111";
		Trees_din <= x"00172961";
		wait for Clk_period;
		Addr <=  "00101000111000";
		Trees_din <= x"13fff104";
		wait for Clk_period;
		Addr <=  "00101000111001";
		Trees_din <= x"00092961";
		wait for Clk_period;
		Addr <=  "00101000111010";
		Trees_din <= x"ffd92961";
		wait for Clk_period;
		Addr <=  "00101000111011";
		Trees_din <= x"1d004004";
		wait for Clk_period;
		Addr <=  "00101000111100";
		Trees_din <= x"00372961";
		wait for Clk_period;
		Addr <=  "00101000111101";
		Trees_din <= x"ff832961";
		wait for Clk_period;
		Addr <=  "00101000111110";
		Trees_din <= x"1400e410";
		wait for Clk_period;
		Addr <=  "00101000111111";
		Trees_din <= x"06f5af04";
		wait for Clk_period;
		Addr <=  "00101001000000";
		Trees_din <= x"ff7c2961";
		wait for Clk_period;
		Addr <=  "00101001000001";
		Trees_din <= x"0f008608";
		wait for Clk_period;
		Addr <=  "00101001000010";
		Trees_din <= x"1c003104";
		wait for Clk_period;
		Addr <=  "00101001000011";
		Trees_din <= x"001a2961";
		wait for Clk_period;
		Addr <=  "00101001000100";
		Trees_din <= x"ffcc2961";
		wait for Clk_period;
		Addr <=  "00101001000101";
		Trees_din <= x"00652961";
		wait for Clk_period;
		Addr <=  "00101001000110";
		Trees_din <= x"0002160c";
		wait for Clk_period;
		Addr <=  "00101001000111";
		Trees_din <= x"0103d308";
		wait for Clk_period;
		Addr <=  "00101001001000";
		Trees_din <= x"10fb1d04";
		wait for Clk_period;
		Addr <=  "00101001001001";
		Trees_din <= x"ffdb2961";
		wait for Clk_period;
		Addr <=  "00101001001010";
		Trees_din <= x"00482961";
		wait for Clk_period;
		Addr <=  "00101001001011";
		Trees_din <= x"ff982961";
		wait for Clk_period;
		Addr <=  "00101001001100";
		Trees_din <= x"08005a08";
		wait for Clk_period;
		Addr <=  "00101001001101";
		Trees_din <= x"020b6104";
		wait for Clk_period;
		Addr <=  "00101001001110";
		Trees_din <= x"ffd82961";
		wait for Clk_period;
		Addr <=  "00101001001111";
		Trees_din <= x"005a2961";
		wait for Clk_period;
		Addr <=  "00101001010000";
		Trees_din <= x"05fc1d04";
		wait for Clk_period;
		Addr <=  "00101001010001";
		Trees_din <= x"00892961";
		wait for Clk_period;
		Addr <=  "00101001010010";
		Trees_din <= x"001c2961";
		wait for Clk_period;
		Addr <=  "00101001010011";
		Trees_din <= x"1c003c08";
		wait for Clk_period;
		Addr <=  "00101001010100";
		Trees_din <= x"1300b404";
		wait for Clk_period;
		Addr <=  "00101001010101";
		Trees_din <= x"ffe92961";
		wait for Clk_period;
		Addr <=  "00101001010110";
		Trees_din <= x"ff942961";
		wait for Clk_period;
		Addr <=  "00101001010111";
		Trees_din <= x"00192961";
		wait for Clk_period;
		Addr <=  "00101001011000";
		Trees_din <= x"02083238";
		wait for Clk_period;
		Addr <=  "00101001011001";
		Trees_din <= x"0c03d72c";
		wait for Clk_period;
		Addr <=  "00101001011010";
		Trees_din <= x"010f7420";
		wait for Clk_period;
		Addr <=  "00101001011011";
		Trees_din <= x"0d034d10";
		wait for Clk_period;
		Addr <=  "00101001011100";
		Trees_din <= x"0d02e908";
		wait for Clk_period;
		Addr <=  "00101001011101";
		Trees_din <= x"03fa6904";
		wait for Clk_period;
		Addr <=  "00101001011110";
		Trees_din <= x"ffcb2a5d";
		wait for Clk_period;
		Addr <=  "00101001011111";
		Trees_din <= x"000a2a5d";
		wait for Clk_period;
		Addr <=  "00101001100000";
		Trees_din <= x"0202c504";
		wait for Clk_period;
		Addr <=  "00101001100001";
		Trees_din <= x"00772a5d";
		wait for Clk_period;
		Addr <=  "00101001100010";
		Trees_din <= x"00002a5d";
		wait for Clk_period;
		Addr <=  "00101001100011";
		Trees_din <= x"07005b08";
		wait for Clk_period;
		Addr <=  "00101001100100";
		Trees_din <= x"00063404";
		wait for Clk_period;
		Addr <=  "00101001100101";
		Trees_din <= x"fff52a5d";
		wait for Clk_period;
		Addr <=  "00101001100110";
		Trees_din <= x"ff712a5d";
		wait for Clk_period;
		Addr <=  "00101001100111";
		Trees_din <= x"01081404";
		wait for Clk_period;
		Addr <=  "00101001101000";
		Trees_din <= x"008c2a5d";
		wait for Clk_period;
		Addr <=  "00101001101001";
		Trees_din <= x"ffd12a5d";
		wait for Clk_period;
		Addr <=  "00101001101010";
		Trees_din <= x"05fb6b08";
		wait for Clk_period;
		Addr <=  "00101001101011";
		Trees_din <= x"11046804";
		wait for Clk_period;
		Addr <=  "00101001101100";
		Trees_din <= x"ff7c2a5d";
		wait for Clk_period;
		Addr <=  "00101001101101";
		Trees_din <= x"002e2a5d";
		wait for Clk_period;
		Addr <=  "00101001101110";
		Trees_din <= x"00492a5d";
		wait for Clk_period;
		Addr <=  "00101001101111";
		Trees_din <= x"0d036b08";
		wait for Clk_period;
		Addr <=  "00101001110000";
		Trees_din <= x"0effcc04";
		wait for Clk_period;
		Addr <=  "00101001110001";
		Trees_din <= x"fffb2a5d";
		wait for Clk_period;
		Addr <=  "00101001110010";
		Trees_din <= x"ff852a5d";
		wait for Clk_period;
		Addr <=  "00101001110011";
		Trees_din <= x"00062a5d";
		wait for Clk_period;
		Addr <=  "00101001110100";
		Trees_din <= x"1202592c";
		wait for Clk_period;
		Addr <=  "00101001110101";
		Trees_din <= x"04ff761c";
		wait for Clk_period;
		Addr <=  "00101001110110";
		Trees_din <= x"03fc5310";
		wait for Clk_period;
		Addr <=  "00101001110111";
		Trees_din <= x"19009608";
		wait for Clk_period;
		Addr <=  "00101001111000";
		Trees_din <= x"18004304";
		wait for Clk_period;
		Addr <=  "00101001111001";
		Trees_din <= x"ff8f2a5d";
		wait for Clk_period;
		Addr <=  "00101001111010";
		Trees_din <= x"001f2a5d";
		wait for Clk_period;
		Addr <=  "00101001111011";
		Trees_din <= x"09004c04";
		wait for Clk_period;
		Addr <=  "00101001111100";
		Trees_din <= x"ffe42a5d";
		wait for Clk_period;
		Addr <=  "00101001111101";
		Trees_din <= x"00502a5d";
		wait for Clk_period;
		Addr <=  "00101001111110";
		Trees_din <= x"0003e504";
		wait for Clk_period;
		Addr <=  "00101001111111";
		Trees_din <= x"00432a5d";
		wait for Clk_period;
		Addr <=  "00101010000000";
		Trees_din <= x"0801f404";
		wait for Clk_period;
		Addr <=  "00101010000001";
		Trees_din <= x"ff952a5d";
		wait for Clk_period;
		Addr <=  "00101010000010";
		Trees_din <= x"00532a5d";
		wait for Clk_period;
		Addr <=  "00101010000011";
		Trees_din <= x"1702f908";
		wait for Clk_period;
		Addr <=  "00101010000100";
		Trees_din <= x"12fe6c04";
		wait for Clk_period;
		Addr <=  "00101010000101";
		Trees_din <= x"001c2a5d";
		wait for Clk_period;
		Addr <=  "00101010000110";
		Trees_din <= x"008e2a5d";
		wait for Clk_period;
		Addr <=  "00101010000111";
		Trees_din <= x"06f2e404";
		wait for Clk_period;
		Addr <=  "00101010001000";
		Trees_din <= x"ffc72a5d";
		wait for Clk_period;
		Addr <=  "00101010001001";
		Trees_din <= x"004c2a5d";
		wait for Clk_period;
		Addr <=  "00101010001010";
		Trees_din <= x"020f9618";
		wait for Clk_period;
		Addr <=  "00101010001011";
		Trees_din <= x"1700b70c";
		wait for Clk_period;
		Addr <=  "00101010001100";
		Trees_din <= x"03fce708";
		wait for Clk_period;
		Addr <=  "00101010001101";
		Trees_din <= x"09005504";
		wait for Clk_period;
		Addr <=  "00101010001110";
		Trees_din <= x"00212a5d";
		wait for Clk_period;
		Addr <=  "00101010001111";
		Trees_din <= x"ffb02a5d";
		wait for Clk_period;
		Addr <=  "00101010010000";
		Trees_din <= x"00712a5d";
		wait for Clk_period;
		Addr <=  "00101010010001";
		Trees_din <= x"09004e04";
		wait for Clk_period;
		Addr <=  "00101010010010";
		Trees_din <= x"001f2a5d";
		wait for Clk_period;
		Addr <=  "00101010010011";
		Trees_din <= x"1d003f04";
		wait for Clk_period;
		Addr <=  "00101010010100";
		Trees_din <= x"ffec2a5d";
		wait for Clk_period;
		Addr <=  "00101010010101";
		Trees_din <= x"ff6b2a5d";
		wait for Clk_period;
		Addr <=  "00101010010110";
		Trees_din <= x"00672a5d";
		wait for Clk_period;
		Addr <=  "00101010010111";
		Trees_din <= x"020baf44";
		wait for Clk_period;
		Addr <=  "00101010011000";
		Trees_din <= x"03f44a08";
		wait for Clk_period;
		Addr <=  "00101010011001";
		Trees_din <= x"08022704";
		wait for Clk_period;
		Addr <=  "00101010011010";
		Trees_din <= x"ff8c2b49";
		wait for Clk_period;
		Addr <=  "00101010011011";
		Trees_din <= x"ffff2b49";
		wait for Clk_period;
		Addr <=  "00101010011100";
		Trees_din <= x"0800151c";
		wait for Clk_period;
		Addr <=  "00101010011101";
		Trees_din <= x"06f7d00c";
		wait for Clk_period;
		Addr <=  "00101010011110";
		Trees_din <= x"1a00f608";
		wait for Clk_period;
		Addr <=  "00101010011111";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00101010100000";
		Trees_din <= x"ff912b49";
		wait for Clk_period;
		Addr <=  "00101010100001";
		Trees_din <= x"ffe52b49";
		wait for Clk_period;
		Addr <=  "00101010100010";
		Trees_din <= x"00432b49";
		wait for Clk_period;
		Addr <=  "00101010100011";
		Trees_din <= x"0afb0708";
		wait for Clk_period;
		Addr <=  "00101010100100";
		Trees_din <= x"0f015904";
		wait for Clk_period;
		Addr <=  "00101010100101";
		Trees_din <= x"fffd2b49";
		wait for Clk_period;
		Addr <=  "00101010100110";
		Trees_din <= x"007b2b49";
		wait for Clk_period;
		Addr <=  "00101010100111";
		Trees_din <= x"1b004904";
		wait for Clk_period;
		Addr <=  "00101010101000";
		Trees_din <= x"ffb32b49";
		wait for Clk_period;
		Addr <=  "00101010101001";
		Trees_din <= x"00222b49";
		wait for Clk_period;
		Addr <=  "00101010101010";
		Trees_din <= x"05fba710";
		wait for Clk_period;
		Addr <=  "00101010101011";
		Trees_din <= x"0e009908";
		wait for Clk_period;
		Addr <=  "00101010101100";
		Trees_din <= x"0efe0804";
		wait for Clk_period;
		Addr <=  "00101010101101";
		Trees_din <= x"00192b49";
		wait for Clk_period;
		Addr <=  "00101010101110";
		Trees_din <= x"ffc12b49";
		wait for Clk_period;
		Addr <=  "00101010101111";
		Trees_din <= x"05fa5804";
		wait for Clk_period;
		Addr <=  "00101010110000";
		Trees_din <= x"00042b49";
		wait for Clk_period;
		Addr <=  "00101010110001";
		Trees_din <= x"004c2b49";
		wait for Clk_period;
		Addr <=  "00101010110010";
		Trees_din <= x"0af7c008";
		wait for Clk_period;
		Addr <=  "00101010110011";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00101010110100";
		Trees_din <= x"ffeb2b49";
		wait for Clk_period;
		Addr <=  "00101010110101";
		Trees_din <= x"ff842b49";
		wait for Clk_period;
		Addr <=  "00101010110110";
		Trees_din <= x"12021b04";
		wait for Clk_period;
		Addr <=  "00101010110111";
		Trees_din <= x"000d2b49";
		wait for Clk_period;
		Addr <=  "00101010111000";
		Trees_din <= x"ffdc2b49";
		wait for Clk_period;
		Addr <=  "00101010111001";
		Trees_din <= x"0001c404";
		wait for Clk_period;
		Addr <=  "00101010111010";
		Trees_din <= x"00732b49";
		wait for Clk_period;
		Addr <=  "00101010111011";
		Trees_din <= x"04f81514";
		wait for Clk_period;
		Addr <=  "00101010111100";
		Trees_din <= x"13ff980c";
		wait for Clk_period;
		Addr <=  "00101010111101";
		Trees_din <= x"0b03b104";
		wait for Clk_period;
		Addr <=  "00101010111110";
		Trees_din <= x"ffc92b49";
		wait for Clk_period;
		Addr <=  "00101010111111";
		Trees_din <= x"0c01bf04";
		wait for Clk_period;
		Addr <=  "00101011000000";
		Trees_din <= x"001a2b49";
		wait for Clk_period;
		Addr <=  "00101011000001";
		Trees_din <= x"005e2b49";
		wait for Clk_period;
		Addr <=  "00101011000010";
		Trees_din <= x"13015504";
		wait for Clk_period;
		Addr <=  "00101011000011";
		Trees_din <= x"00812b49";
		wait for Clk_period;
		Addr <=  "00101011000100";
		Trees_din <= x"001c2b49";
		wait for Clk_period;
		Addr <=  "00101011000101";
		Trees_din <= x"1601120c";
		wait for Clk_period;
		Addr <=  "00101011000110";
		Trees_din <= x"13fd9808";
		wait for Clk_period;
		Addr <=  "00101011000111";
		Trees_din <= x"1a00c304";
		wait for Clk_period;
		Addr <=  "00101011001000";
		Trees_din <= x"ffac2b49";
		wait for Clk_period;
		Addr <=  "00101011001001";
		Trees_din <= x"00222b49";
		wait for Clk_period;
		Addr <=  "00101011001010";
		Trees_din <= x"00782b49";
		wait for Clk_period;
		Addr <=  "00101011001011";
		Trees_din <= x"12015b08";
		wait for Clk_period;
		Addr <=  "00101011001100";
		Trees_din <= x"00108804";
		wait for Clk_period;
		Addr <=  "00101011001101";
		Trees_din <= x"003f2b49";
		wait for Clk_period;
		Addr <=  "00101011001110";
		Trees_din <= x"ffa62b49";
		wait for Clk_period;
		Addr <=  "00101011001111";
		Trees_din <= x"10fab704";
		wait for Clk_period;
		Addr <=  "00101011010000";
		Trees_din <= x"00302b49";
		wait for Clk_period;
		Addr <=  "00101011010001";
		Trees_din <= x"ff972b49";
		wait for Clk_period;
		Addr <=  "00101011010010";
		Trees_din <= x"0204753c";
		wait for Clk_period;
		Addr <=  "00101011010011";
		Trees_din <= x"02040934";
		wait for Clk_period;
		Addr <=  "00101011010100";
		Trees_din <= x"0d03371c";
		wait for Clk_period;
		Addr <=  "00101011010101";
		Trees_din <= x"0d02e910";
		wait for Clk_period;
		Addr <=  "00101011010110";
		Trees_din <= x"0203a108";
		wait for Clk_period;
		Addr <=  "00101011010111";
		Trees_din <= x"1203f704";
		wait for Clk_period;
		Addr <=  "00101011011000";
		Trees_din <= x"ffdd2c25";
		wait for Clk_period;
		Addr <=  "00101011011001";
		Trees_din <= x"00482c25";
		wait for Clk_period;
		Addr <=  "00101011011010";
		Trees_din <= x"0d016504";
		wait for Clk_period;
		Addr <=  "00101011011011";
		Trees_din <= x"007b2c25";
		wait for Clk_period;
		Addr <=  "00101011011100";
		Trees_din <= x"ffc62c25";
		wait for Clk_period;
		Addr <=  "00101011011101";
		Trees_din <= x"16039608";
		wait for Clk_period;
		Addr <=  "00101011011110";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00101011011111";
		Trees_din <= x"00902c25";
		wait for Clk_period;
		Addr <=  "00101011100000";
		Trees_din <= x"002a2c25";
		wait for Clk_period;
		Addr <=  "00101011100001";
		Trees_din <= x"ffc32c25";
		wait for Clk_period;
		Addr <=  "00101011100010";
		Trees_din <= x"1700f10c";
		wait for Clk_period;
		Addr <=  "00101011100011";
		Trees_din <= x"0c038c04";
		wait for Clk_period;
		Addr <=  "00101011100100";
		Trees_din <= x"ff882c25";
		wait for Clk_period;
		Addr <=  "00101011100101";
		Trees_din <= x"11022704";
		wait for Clk_period;
		Addr <=  "00101011100110";
		Trees_din <= x"00132c25";
		wait for Clk_period;
		Addr <=  "00101011100111";
		Trees_din <= x"ffe22c25";
		wait for Clk_period;
		Addr <=  "00101011101000";
		Trees_din <= x"10046a04";
		wait for Clk_period;
		Addr <=  "00101011101001";
		Trees_din <= x"ffab2c25";
		wait for Clk_period;
		Addr <=  "00101011101010";
		Trees_din <= x"0bf95804";
		wait for Clk_period;
		Addr <=  "00101011101011";
		Trees_din <= x"00632c25";
		wait for Clk_period;
		Addr <=  "00101011101100";
		Trees_din <= x"000b2c25";
		wait for Clk_period;
		Addr <=  "00101011101101";
		Trees_din <= x"1c004004";
		wait for Clk_period;
		Addr <=  "00101011101110";
		Trees_din <= x"ff8d2c25";
		wait for Clk_period;
		Addr <=  "00101011101111";
		Trees_din <= x"ffef2c25";
		wait for Clk_period;
		Addr <=  "00101011110000";
		Trees_din <= x"0e041128";
		wait for Clk_period;
		Addr <=  "00101011110001";
		Trees_din <= x"00fe7b0c";
		wait for Clk_period;
		Addr <=  "00101011110010";
		Trees_din <= x"13f9d204";
		wait for Clk_period;
		Addr <=  "00101011110011";
		Trees_din <= x"ffed2c25";
		wait for Clk_period;
		Addr <=  "00101011110100";
		Trees_din <= x"07005404";
		wait for Clk_period;
		Addr <=  "00101011110101";
		Trees_din <= x"001c2c25";
		wait for Clk_period;
		Addr <=  "00101011110110";
		Trees_din <= x"006e2c25";
		wait for Clk_period;
		Addr <=  "00101011110111";
		Trees_din <= x"11044410";
		wait for Clk_period;
		Addr <=  "00101011111000";
		Trees_din <= x"0e025a08";
		wait for Clk_period;
		Addr <=  "00101011111001";
		Trees_din <= x"11030f04";
		wait for Clk_period;
		Addr <=  "00101011111010";
		Trees_din <= x"00082c25";
		wait for Clk_period;
		Addr <=  "00101011111011";
		Trees_din <= x"00732c25";
		wait for Clk_period;
		Addr <=  "00101011111100";
		Trees_din <= x"13ff8804";
		wait for Clk_period;
		Addr <=  "00101011111101";
		Trees_din <= x"ff932c25";
		wait for Clk_period;
		Addr <=  "00101011111110";
		Trees_din <= x"fff82c25";
		wait for Clk_period;
		Addr <=  "00101011111111";
		Trees_din <= x"03f5be04";
		wait for Clk_period;
		Addr <=  "00101100000000";
		Trees_din <= x"ffbf2c25";
		wait for Clk_period;
		Addr <=  "00101100000001";
		Trees_din <= x"09005604";
		wait for Clk_period;
		Addr <=  "00101100000010";
		Trees_din <= x"00712c25";
		wait for Clk_period;
		Addr <=  "00101100000011";
		Trees_din <= x"ffec2c25";
		wait for Clk_period;
		Addr <=  "00101100000100";
		Trees_din <= x"10fade04";
		wait for Clk_period;
		Addr <=  "00101100000101";
		Trees_din <= x"002a2c25";
		wait for Clk_period;
		Addr <=  "00101100000110";
		Trees_din <= x"0103d304";
		wait for Clk_period;
		Addr <=  "00101100000111";
		Trees_din <= x"00092c25";
		wait for Clk_period;
		Addr <=  "00101100001000";
		Trees_din <= x"ff8d2c25";
		wait for Clk_period;
		Addr <=  "00101100001001";
		Trees_din <= x"020baf3c";
		wait for Clk_period;
		Addr <=  "00101100001010";
		Trees_din <= x"03f44a08";
		wait for Clk_period;
		Addr <=  "00101100001011";
		Trees_din <= x"0801f404";
		wait for Clk_period;
		Addr <=  "00101100001100";
		Trees_din <= x"ff932cf9";
		wait for Clk_period;
		Addr <=  "00101100001101";
		Trees_din <= x"fffd2cf9";
		wait for Clk_period;
		Addr <=  "00101100001110";
		Trees_din <= x"0d000514";
		wait for Clk_period;
		Addr <=  "00101100001111";
		Trees_din <= x"20040008";
		wait for Clk_period;
		Addr <=  "00101100010000";
		Trees_din <= x"0103ae04";
		wait for Clk_period;
		Addr <=  "00101100010001";
		Trees_din <= x"002d2cf9";
		wait for Clk_period;
		Addr <=  "00101100010010";
		Trees_din <= x"ff9e2cf9";
		wait for Clk_period;
		Addr <=  "00101100010011";
		Trees_din <= x"02037004";
		wait for Clk_period;
		Addr <=  "00101100010100";
		Trees_din <= x"fffd2cf9";
		wait for Clk_period;
		Addr <=  "00101100010101";
		Trees_din <= x"0007fa04";
		wait for Clk_period;
		Addr <=  "00101100010110";
		Trees_din <= x"000b2cf9";
		wait for Clk_period;
		Addr <=  "00101100010111";
		Trees_din <= x"009e2cf9";
		wait for Clk_period;
		Addr <=  "00101100011000";
		Trees_din <= x"0d003410";
		wait for Clk_period;
		Addr <=  "00101100011001";
		Trees_din <= x"11028808";
		wait for Clk_period;
		Addr <=  "00101100011010";
		Trees_din <= x"08006404";
		wait for Clk_period;
		Addr <=  "00101100011011";
		Trees_din <= x"00072cf9";
		wait for Clk_period;
		Addr <=  "00101100011100";
		Trees_din <= x"ff7e2cf9";
		wait for Clk_period;
		Addr <=  "00101100011101";
		Trees_din <= x"1102b304";
		wait for Clk_period;
		Addr <=  "00101100011110";
		Trees_din <= x"00712cf9";
		wait for Clk_period;
		Addr <=  "00101100011111";
		Trees_din <= x"ffdd2cf9";
		wait for Clk_period;
		Addr <=  "00101100100000";
		Trees_din <= x"05fba708";
		wait for Clk_period;
		Addr <=  "00101100100001";
		Trees_din <= x"05f5f504";
		wait for Clk_period;
		Addr <=  "00101100100010";
		Trees_din <= x"ffb42cf9";
		wait for Clk_period;
		Addr <=  "00101100100011";
		Trees_din <= x"00132cf9";
		wait for Clk_period;
		Addr <=  "00101100100100";
		Trees_din <= x"12fe4404";
		wait for Clk_period;
		Addr <=  "00101100100101";
		Trees_din <= x"002d2cf9";
		wait for Clk_period;
		Addr <=  "00101100100110";
		Trees_din <= x"ffe62cf9";
		wait for Clk_period;
		Addr <=  "00101100100111";
		Trees_din <= x"0001c404";
		wait for Clk_period;
		Addr <=  "00101100101000";
		Trees_din <= x"006e2cf9";
		wait for Clk_period;
		Addr <=  "00101100101001";
		Trees_din <= x"04f81510";
		wait for Clk_period;
		Addr <=  "00101100101010";
		Trees_din <= x"1005890c";
		wait for Clk_period;
		Addr <=  "00101100101011";
		Trees_din <= x"12008804";
		wait for Clk_period;
		Addr <=  "00101100101100";
		Trees_din <= x"00002cf9";
		wait for Clk_period;
		Addr <=  "00101100101101";
		Trees_din <= x"17002704";
		wait for Clk_period;
		Addr <=  "00101100101110";
		Trees_din <= x"001e2cf9";
		wait for Clk_period;
		Addr <=  "00101100101111";
		Trees_din <= x"00722cf9";
		wait for Clk_period;
		Addr <=  "00101100110000";
		Trees_din <= x"fffc2cf9";
		wait for Clk_period;
		Addr <=  "00101100110001";
		Trees_din <= x"12015b0c";
		wait for Clk_period;
		Addr <=  "00101100110010";
		Trees_din <= x"00115708";
		wait for Clk_period;
		Addr <=  "00101100110011";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00101100110100";
		Trees_din <= x"ffd52cf9";
		wait for Clk_period;
		Addr <=  "00101100110101";
		Trees_din <= x"005c2cf9";
		wait for Clk_period;
		Addr <=  "00101100110110";
		Trees_din <= x"ffb02cf9";
		wait for Clk_period;
		Addr <=  "00101100110111";
		Trees_din <= x"0f022d08";
		wait for Clk_period;
		Addr <=  "00101100111000";
		Trees_din <= x"10fac504";
		wait for Clk_period;
		Addr <=  "00101100111001";
		Trees_din <= x"002b2cf9";
		wait for Clk_period;
		Addr <=  "00101100111010";
		Trees_din <= x"ff9c2cf9";
		wait for Clk_period;
		Addr <=  "00101100111011";
		Trees_din <= x"000ceb04";
		wait for Clk_period;
		Addr <=  "00101100111100";
		Trees_din <= x"00642cf9";
		wait for Clk_period;
		Addr <=  "00101100111101";
		Trees_din <= x"ffd52cf9";
		wait for Clk_period;
		Addr <=  "00101100111110";
		Trees_din <= x"02083240";
		wait for Clk_period;
		Addr <=  "00101100111111";
		Trees_din <= x"0b056f34";
		wait for Clk_period;
		Addr <=  "00101101000000";
		Trees_din <= x"1b002e14";
		wait for Clk_period;
		Addr <=  "00101101000001";
		Trees_din <= x"0201e304";
		wait for Clk_period;
		Addr <=  "00101101000010";
		Trees_din <= x"ff872dcd";
		wait for Clk_period;
		Addr <=  "00101101000011";
		Trees_din <= x"02036308";
		wait for Clk_period;
		Addr <=  "00101101000100";
		Trees_din <= x"06f59f04";
		wait for Clk_period;
		Addr <=  "00101101000101";
		Trees_din <= x"ffdb2dcd";
		wait for Clk_period;
		Addr <=  "00101101000110";
		Trees_din <= x"00592dcd";
		wait for Clk_period;
		Addr <=  "00101101000111";
		Trees_din <= x"0d01d504";
		wait for Clk_period;
		Addr <=  "00101101001000";
		Trees_din <= x"000c2dcd";
		wait for Clk_period;
		Addr <=  "00101101001001";
		Trees_din <= x"ff9a2dcd";
		wait for Clk_period;
		Addr <=  "00101101001010";
		Trees_din <= x"08001510";
		wait for Clk_period;
		Addr <=  "00101101001011";
		Trees_din <= x"06f7d008";
		wait for Clk_period;
		Addr <=  "00101101001100";
		Trees_din <= x"05fd2704";
		wait for Clk_period;
		Addr <=  "00101101001101";
		Trees_din <= x"ff9a2dcd";
		wait for Clk_period;
		Addr <=  "00101101001110";
		Trees_din <= x"00082dcd";
		wait for Clk_period;
		Addr <=  "00101101001111";
		Trees_din <= x"03fda804";
		wait for Clk_period;
		Addr <=  "00101101010000";
		Trees_din <= x"ffcb2dcd";
		wait for Clk_period;
		Addr <=  "00101101010001";
		Trees_din <= x"003d2dcd";
		wait for Clk_period;
		Addr <=  "00101101010010";
		Trees_din <= x"1c003208";
		wait for Clk_period;
		Addr <=  "00101101010011";
		Trees_din <= x"0d036504";
		wait for Clk_period;
		Addr <=  "00101101010100";
		Trees_din <= x"00302dcd";
		wait for Clk_period;
		Addr <=  "00101101010101";
		Trees_din <= x"ffa32dcd";
		wait for Clk_period;
		Addr <=  "00101101010110";
		Trees_din <= x"1b004504";
		wait for Clk_period;
		Addr <=  "00101101010111";
		Trees_din <= x"ffec2dcd";
		wait for Clk_period;
		Addr <=  "00101101011000";
		Trees_din <= x"00392dcd";
		wait for Clk_period;
		Addr <=  "00101101011001";
		Trees_din <= x"12fdf608";
		wait for Clk_period;
		Addr <=  "00101101011010";
		Trees_din <= x"12fda004";
		wait for Clk_period;
		Addr <=  "00101101011011";
		Trees_din <= x"ffd52dcd";
		wait for Clk_period;
		Addr <=  "00101101011100";
		Trees_din <= x"00572dcd";
		wait for Clk_period;
		Addr <=  "00101101011101";
		Trees_din <= x"ff8e2dcd";
		wait for Clk_period;
		Addr <=  "00101101011110";
		Trees_din <= x"08000508";
		wait for Clk_period;
		Addr <=  "00101101011111";
		Trees_din <= x"15008004";
		wait for Clk_period;
		Addr <=  "00101101100000";
		Trees_din <= x"00022dcd";
		wait for Clk_period;
		Addr <=  "00101101100001";
		Trees_din <= x"00692dcd";
		wait for Clk_period;
		Addr <=  "00101101100010";
		Trees_din <= x"10068320";
		wait for Clk_period;
		Addr <=  "00101101100011";
		Trees_din <= x"06f34c10";
		wait for Clk_period;
		Addr <=  "00101101100100";
		Trees_din <= x"0d01f208";
		wait for Clk_period;
		Addr <=  "00101101100101";
		Trees_din <= x"05fc5d04";
		wait for Clk_period;
		Addr <=  "00101101100110";
		Trees_din <= x"ffb22dcd";
		wait for Clk_period;
		Addr <=  "00101101100111";
		Trees_din <= x"00342dcd";
		wait for Clk_period;
		Addr <=  "00101101101000";
		Trees_din <= x"000e0e04";
		wait for Clk_period;
		Addr <=  "00101101101001";
		Trees_din <= x"00362dcd";
		wait for Clk_period;
		Addr <=  "00101101101010";
		Trees_din <= x"ffa62dcd";
		wait for Clk_period;
		Addr <=  "00101101101011";
		Trees_din <= x"0801f408";
		wait for Clk_period;
		Addr <=  "00101101101100";
		Trees_din <= x"000d6304";
		wait for Clk_period;
		Addr <=  "00101101101101";
		Trees_din <= x"001b2dcd";
		wait for Clk_period;
		Addr <=  "00101101101110";
		Trees_din <= x"ffd92dcd";
		wait for Clk_period;
		Addr <=  "00101101101111";
		Trees_din <= x"1b003204";
		wait for Clk_period;
		Addr <=  "00101101110000";
		Trees_din <= x"000a2dcd";
		wait for Clk_period;
		Addr <=  "00101101110001";
		Trees_din <= x"00712dcd";
		wait for Clk_period;
		Addr <=  "00101101110010";
		Trees_din <= x"00632dcd";
		wait for Clk_period;
		Addr <=  "00101101110011";
		Trees_din <= x"21000158";
		wait for Clk_period;
		Addr <=  "00101101110100";
		Trees_din <= x"02058f30";
		wait for Clk_period;
		Addr <=  "00101101110101";
		Trees_din <= x"07005918";
		wait for Clk_period;
		Addr <=  "00101101110110";
		Trees_din <= x"10063110";
		wait for Clk_period;
		Addr <=  "00101101110111";
		Trees_din <= x"04fb2808";
		wait for Clk_period;
		Addr <=  "00101101111000";
		Trees_din <= x"13ffb904";
		wait for Clk_period;
		Addr <=  "00101101111001";
		Trees_din <= x"ffa92e91";
		wait for Clk_period;
		Addr <=  "00101101111010";
		Trees_din <= x"001c2e91";
		wait for Clk_period;
		Addr <=  "00101101111011";
		Trees_din <= x"0204e504";
		wait for Clk_period;
		Addr <=  "00101101111100";
		Trees_din <= x"00012e91";
		wait for Clk_period;
		Addr <=  "00101101111101";
		Trees_din <= x"004a2e91";
		wait for Clk_period;
		Addr <=  "00101101111110";
		Trees_din <= x"0bfa9f04";
		wait for Clk_period;
		Addr <=  "00101101111111";
		Trees_din <= x"ffe32e91";
		wait for Clk_period;
		Addr <=  "00101110000000";
		Trees_din <= x"ff962e91";
		wait for Clk_period;
		Addr <=  "00101110000001";
		Trees_din <= x"05fc3808";
		wait for Clk_period;
		Addr <=  "00101110000010";
		Trees_din <= x"09005904";
		wait for Clk_period;
		Addr <=  "00101110000011";
		Trees_din <= x"ff802e91";
		wait for Clk_period;
		Addr <=  "00101110000100";
		Trees_din <= x"fff32e91";
		wait for Clk_period;
		Addr <=  "00101110000101";
		Trees_din <= x"13ff9508";
		wait for Clk_period;
		Addr <=  "00101110000110";
		Trees_din <= x"03fe8b04";
		wait for Clk_period;
		Addr <=  "00101110000111";
		Trees_din <= x"ffcd2e91";
		wait for Clk_period;
		Addr <=  "00101110001000";
		Trees_din <= x"00582e91";
		wait for Clk_period;
		Addr <=  "00101110001001";
		Trees_din <= x"1b004704";
		wait for Clk_period;
		Addr <=  "00101110001010";
		Trees_din <= x"ff932e91";
		wait for Clk_period;
		Addr <=  "00101110001011";
		Trees_din <= x"00232e91";
		wait for Clk_period;
		Addr <=  "00101110001100";
		Trees_din <= x"10068320";
		wait for Clk_period;
		Addr <=  "00101110001101";
		Trees_din <= x"07005910";
		wait for Clk_period;
		Addr <=  "00101110001110";
		Trees_din <= x"09005508";
		wait for Clk_period;
		Addr <=  "00101110001111";
		Trees_din <= x"02079804";
		wait for Clk_period;
		Addr <=  "00101110010000";
		Trees_din <= x"ffde2e91";
		wait for Clk_period;
		Addr <=  "00101110010001";
		Trees_din <= x"001e2e91";
		wait for Clk_period;
		Addr <=  "00101110010010";
		Trees_din <= x"09005704";
		wait for Clk_period;
		Addr <=  "00101110010011";
		Trees_din <= x"ffb12e91";
		wait for Clk_period;
		Addr <=  "00101110010100";
		Trees_din <= x"00002e91";
		wait for Clk_period;
		Addr <=  "00101110010101";
		Trees_din <= x"1d004608";
		wait for Clk_period;
		Addr <=  "00101110010110";
		Trees_din <= x"1e007004";
		wait for Clk_period;
		Addr <=  "00101110010111";
		Trees_din <= x"00602e91";
		wait for Clk_period;
		Addr <=  "00101110011000";
		Trees_din <= x"ffcc2e91";
		wait for Clk_period;
		Addr <=  "00101110011001";
		Trees_din <= x"1e006c04";
		wait for Clk_period;
		Addr <=  "00101110011010";
		Trees_din <= x"ff872e91";
		wait for Clk_period;
		Addr <=  "00101110011011";
		Trees_din <= x"000f2e91";
		wait for Clk_period;
		Addr <=  "00101110011100";
		Trees_din <= x"19009404";
		wait for Clk_period;
		Addr <=  "00101110011101";
		Trees_din <= x"001f2e91";
		wait for Clk_period;
		Addr <=  "00101110011110";
		Trees_din <= x"006f2e91";
		wait for Clk_period;
		Addr <=  "00101110011111";
		Trees_din <= x"01076004";
		wait for Clk_period;
		Addr <=  "00101110100000";
		Trees_din <= x"ffcd2e91";
		wait for Clk_period;
		Addr <=  "00101110100001";
		Trees_din <= x"010d4f04";
		wait for Clk_period;
		Addr <=  "00101110100010";
		Trees_din <= x"007a2e91";
		wait for Clk_period;
		Addr <=  "00101110100011";
		Trees_din <= x"00142e91";
		wait for Clk_period;
		Addr <=  "00101110100100";
		Trees_din <= x"21000154";
		wait for Clk_period;
		Addr <=  "00101110100101";
		Trees_din <= x"02058f30";
		wait for Clk_period;
		Addr <=  "00101110100110";
		Trees_din <= x"03fa5a14";
		wait for Clk_period;
		Addr <=  "00101110100111";
		Trees_din <= x"0c028d08";
		wait for Clk_period;
		Addr <=  "00101110101000";
		Trees_din <= x"00161e04";
		wait for Clk_period;
		Addr <=  "00101110101001";
		Trees_din <= x"ff7c2f4d";
		wait for Clk_period;
		Addr <=  "00101110101010";
		Trees_din <= x"00012f4d";
		wait for Clk_period;
		Addr <=  "00101110101011";
		Trees_din <= x"13fe4d08";
		wait for Clk_period;
		Addr <=  "00101110101100";
		Trees_din <= x"06f4ea04";
		wait for Clk_period;
		Addr <=  "00101110101101";
		Trees_din <= x"00872f4d";
		wait for Clk_period;
		Addr <=  "00101110101110";
		Trees_din <= x"000f2f4d";
		wait for Clk_period;
		Addr <=  "00101110101111";
		Trees_din <= x"ff912f4d";
		wait for Clk_period;
		Addr <=  "00101110110000";
		Trees_din <= x"03fafe0c";
		wait for Clk_period;
		Addr <=  "00101110110001";
		Trees_din <= x"13016508";
		wait for Clk_period;
		Addr <=  "00101110110010";
		Trees_din <= x"05fde504";
		wait for Clk_period;
		Addr <=  "00101110110011";
		Trees_din <= x"ffaa2f4d";
		wait for Clk_period;
		Addr <=  "00101110110100";
		Trees_din <= x"005d2f4d";
		wait for Clk_period;
		Addr <=  "00101110110101";
		Trees_din <= x"00892f4d";
		wait for Clk_period;
		Addr <=  "00101110110110";
		Trees_din <= x"07005908";
		wait for Clk_period;
		Addr <=  "00101110110111";
		Trees_din <= x"1a00a604";
		wait for Clk_period;
		Addr <=  "00101110111000";
		Trees_din <= x"00372f4d";
		wait for Clk_period;
		Addr <=  "00101110111001";
		Trees_din <= x"fff72f4d";
		wait for Clk_period;
		Addr <=  "00101110111010";
		Trees_din <= x"0efcb004";
		wait for Clk_period;
		Addr <=  "00101110111011";
		Trees_din <= x"00292f4d";
		wait for Clk_period;
		Addr <=  "00101110111100";
		Trees_din <= x"ffaf2f4d";
		wait for Clk_period;
		Addr <=  "00101110111101";
		Trees_din <= x"1d003304";
		wait for Clk_period;
		Addr <=  "00101110111110";
		Trees_din <= x"ffa82f4d";
		wait for Clk_period;
		Addr <=  "00101110111111";
		Trees_din <= x"0d011010";
		wait for Clk_period;
		Addr <=  "00101111000000";
		Trees_din <= x"06f35808";
		wait for Clk_period;
		Addr <=  "00101111000001";
		Trees_din <= x"15008904";
		wait for Clk_period;
		Addr <=  "00101111000010";
		Trees_din <= x"ff9e2f4d";
		wait for Clk_period;
		Addr <=  "00101111000011";
		Trees_din <= x"001a2f4d";
		wait for Clk_period;
		Addr <=  "00101111000100";
		Trees_din <= x"03fb3a04";
		wait for Clk_period;
		Addr <=  "00101111000101";
		Trees_din <= x"00152f4d";
		wait for Clk_period;
		Addr <=  "00101111000110";
		Trees_din <= x"00622f4d";
		wait for Clk_period;
		Addr <=  "00101111000111";
		Trees_din <= x"0d017a08";
		wait for Clk_period;
		Addr <=  "00101111001000";
		Trees_din <= x"0c00c704";
		wait for Clk_period;
		Addr <=  "00101111001001";
		Trees_din <= x"002d2f4d";
		wait for Clk_period;
		Addr <=  "00101111001010";
		Trees_din <= x"ff8a2f4d";
		wait for Clk_period;
		Addr <=  "00101111001011";
		Trees_din <= x"09004f04";
		wait for Clk_period;
		Addr <=  "00101111001100";
		Trees_din <= x"ffd42f4d";
		wait for Clk_period;
		Addr <=  "00101111001101";
		Trees_din <= x"00122f4d";
		wait for Clk_period;
		Addr <=  "00101111001110";
		Trees_din <= x"01076004";
		wait for Clk_period;
		Addr <=  "00101111001111";
		Trees_din <= x"ffd22f4d";
		wait for Clk_period;
		Addr <=  "00101111010000";
		Trees_din <= x"010d4f04";
		wait for Clk_period;
		Addr <=  "00101111010001";
		Trees_din <= x"00712f4d";
		wait for Clk_period;
		Addr <=  "00101111010010";
		Trees_din <= x"00122f4d";
		wait for Clk_period;
		Addr <=  "00101111010011";
		Trees_din <= x"020baf34";
		wait for Clk_period;
		Addr <=  "00101111010100";
		Trees_din <= x"03f44a08";
		wait for Clk_period;
		Addr <=  "00101111010101";
		Trees_din <= x"0015c504";
		wait for Clk_period;
		Addr <=  "00101111010110";
		Trees_din <= x"ff9c3019";
		wait for Clk_period;
		Addr <=  "00101111010111";
		Trees_din <= x"ffec3019";
		wait for Clk_period;
		Addr <=  "00101111011000";
		Trees_din <= x"0f000418";
		wait for Clk_period;
		Addr <=  "00101111011001";
		Trees_din <= x"1200c80c";
		wait for Clk_period;
		Addr <=  "00101111011010";
		Trees_din <= x"0b04f208";
		wait for Clk_period;
		Addr <=  "00101111011011";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00101111011100";
		Trees_din <= x"00873019";
		wait for Clk_period;
		Addr <=  "00101111011101";
		Trees_din <= x"00043019";
		wait for Clk_period;
		Addr <=  "00101111011110";
		Trees_din <= x"ffc53019";
		wait for Clk_period;
		Addr <=  "00101111011111";
		Trees_din <= x"0a02ad08";
		wait for Clk_period;
		Addr <=  "00101111100000";
		Trees_din <= x"02058f04";
		wait for Clk_period;
		Addr <=  "00101111100001";
		Trees_din <= x"ffac3019";
		wait for Clk_period;
		Addr <=  "00101111100010";
		Trees_din <= x"00183019";
		wait for Clk_period;
		Addr <=  "00101111100011";
		Trees_din <= x"00463019";
		wait for Clk_period;
		Addr <=  "00101111100100";
		Trees_din <= x"02fda204";
		wait for Clk_period;
		Addr <=  "00101111100101";
		Trees_din <= x"ff993019";
		wait for Clk_period;
		Addr <=  "00101111100110";
		Trees_din <= x"0d000508";
		wait for Clk_period;
		Addr <=  "00101111100111";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00101111101000";
		Trees_din <= x"ffd63019";
		wait for Clk_period;
		Addr <=  "00101111101001";
		Trees_din <= x"00513019";
		wait for Clk_period;
		Addr <=  "00101111101010";
		Trees_din <= x"0c004a04";
		wait for Clk_period;
		Addr <=  "00101111101011";
		Trees_din <= x"ffb43019";
		wait for Clk_period;
		Addr <=  "00101111101100";
		Trees_din <= x"fffc3019";
		wait for Clk_period;
		Addr <=  "00101111101101";
		Trees_din <= x"01025918";
		wait for Clk_period;
		Addr <=  "00101111101110";
		Trees_din <= x"0afc7c0c";
		wait for Clk_period;
		Addr <=  "00101111101111";
		Trees_din <= x"08002d04";
		wait for Clk_period;
		Addr <=  "00101111110000";
		Trees_din <= x"00513019";
		wait for Clk_period;
		Addr <=  "00101111110001";
		Trees_din <= x"19009204";
		wait for Clk_period;
		Addr <=  "00101111110010";
		Trees_din <= x"ffe83019";
		wait for Clk_period;
		Addr <=  "00101111110011";
		Trees_din <= x"ff723019";
		wait for Clk_period;
		Addr <=  "00101111110100";
		Trees_din <= x"00103308";
		wait for Clk_period;
		Addr <=  "00101111110101";
		Trees_din <= x"0801cf04";
		wait for Clk_period;
		Addr <=  "00101111110110";
		Trees_din <= x"00693019";
		wait for Clk_period;
		Addr <=  "00101111110111";
		Trees_din <= x"001b3019";
		wait for Clk_period;
		Addr <=  "00101111111000";
		Trees_din <= x"ffd23019";
		wait for Clk_period;
		Addr <=  "00101111111001";
		Trees_din <= x"0f000004";
		wait for Clk_period;
		Addr <=  "00101111111010";
		Trees_din <= x"ffc03019";
		wait for Clk_period;
		Addr <=  "00101111111011";
		Trees_din <= x"0efb0d08";
		wait for Clk_period;
		Addr <=  "00101111111100";
		Trees_din <= x"15008704";
		wait for Clk_period;
		Addr <=  "00101111111101";
		Trees_din <= x"ff9e3019";
		wait for Clk_period;
		Addr <=  "00101111111110";
		Trees_din <= x"00253019";
		wait for Clk_period;
		Addr <=  "00101111111111";
		Trees_din <= x"0e025a08";
		wait for Clk_period;
		Addr <=  "00110000000000";
		Trees_din <= x"06f00004";
		wait for Clk_period;
		Addr <=  "00110000000001";
		Trees_din <= x"fff03019";
		wait for Clk_period;
		Addr <=  "00110000000010";
		Trees_din <= x"005b3019";
		wait for Clk_period;
		Addr <=  "00110000000011";
		Trees_din <= x"09005004";
		wait for Clk_period;
		Addr <=  "00110000000100";
		Trees_din <= x"ffc23019";
		wait for Clk_period;
		Addr <=  "00110000000101";
		Trees_din <= x"00373019";
		wait for Clk_period;
		Addr <=  "00110000000110";
		Trees_din <= x"00fc3a1c";
		wait for Clk_period;
		Addr <=  "00110000000111";
		Trees_din <= x"00f95808";
		wait for Clk_period;
		Addr <=  "00110000001000";
		Trees_din <= x"02032e04";
		wait for Clk_period;
		Addr <=  "00110000001001";
		Trees_din <= x"ffa630f5";
		wait for Clk_period;
		Addr <=  "00110000001010";
		Trees_din <= x"002330f5";
		wait for Clk_period;
		Addr <=  "00110000001011";
		Trees_din <= x"19009f0c";
		wait for Clk_period;
		Addr <=  "00110000001100";
		Trees_din <= x"1b004308";
		wait for Clk_period;
		Addr <=  "00110000001101";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00110000001110";
		Trees_din <= x"006e30f5";
		wait for Clk_period;
		Addr <=  "00110000001111";
		Trees_din <= x"001f30f5";
		wait for Clk_period;
		Addr <=  "00110000010000";
		Trees_din <= x"fff130f5";
		wait for Clk_period;
		Addr <=  "00110000010001";
		Trees_din <= x"0d01bb04";
		wait for Clk_period;
		Addr <=  "00110000010010";
		Trees_din <= x"001830f5";
		wait for Clk_period;
		Addr <=  "00110000010011";
		Trees_din <= x"ffc730f5";
		wait for Clk_period;
		Addr <=  "00110000010100";
		Trees_din <= x"1500aa30";
		wait for Clk_period;
		Addr <=  "00110000010101";
		Trees_din <= x"1500a71c";
		wait for Clk_period;
		Addr <=  "00110000010110";
		Trees_din <= x"1500a610";
		wait for Clk_period;
		Addr <=  "00110000010111";
		Trees_din <= x"02047508";
		wait for Clk_period;
		Addr <=  "00110000011000";
		Trees_din <= x"0e046904";
		wait for Clk_period;
		Addr <=  "00110000011001";
		Trees_din <= x"ffdd30f5";
		wait for Clk_period;
		Addr <=  "00110000011010";
		Trees_din <= x"004730f5";
		wait for Clk_period;
		Addr <=  "00110000011011";
		Trees_din <= x"05003a04";
		wait for Clk_period;
		Addr <=  "00110000011100";
		Trees_din <= x"ffff30f5";
		wait for Clk_period;
		Addr <=  "00110000011101";
		Trees_din <= x"003a30f5";
		wait for Clk_period;
		Addr <=  "00110000011110";
		Trees_din <= x"0a024104";
		wait for Clk_period;
		Addr <=  "00110000011111";
		Trees_din <= x"ffef30f5";
		wait for Clk_period;
		Addr <=  "00110000100000";
		Trees_din <= x"0c015d04";
		wait for Clk_period;
		Addr <=  "00110000100001";
		Trees_din <= x"007630f5";
		wait for Clk_period;
		Addr <=  "00110000100010";
		Trees_din <= x"002130f5";
		wait for Clk_period;
		Addr <=  "00110000100011";
		Trees_din <= x"0efe2604";
		wait for Clk_period;
		Addr <=  "00110000100100";
		Trees_din <= x"ff8730f5";
		wait for Clk_period;
		Addr <=  "00110000100101";
		Trees_din <= x"0b048208";
		wait for Clk_period;
		Addr <=  "00110000100110";
		Trees_din <= x"02083204";
		wait for Clk_period;
		Addr <=  "00110000100111";
		Trees_din <= x"ffa630f5";
		wait for Clk_period;
		Addr <=  "00110000101000";
		Trees_din <= x"002230f5";
		wait for Clk_period;
		Addr <=  "00110000101001";
		Trees_din <= x"0afc8304";
		wait for Clk_period;
		Addr <=  "00110000101010";
		Trees_din <= x"001830f5";
		wait for Clk_period;
		Addr <=  "00110000101011";
		Trees_din <= x"005b30f5";
		wait for Clk_period;
		Addr <=  "00110000101100";
		Trees_din <= x"1d003b1c";
		wait for Clk_period;
		Addr <=  "00110000101101";
		Trees_din <= x"08009b0c";
		wait for Clk_period;
		Addr <=  "00110000101110";
		Trees_din <= x"06f6ad08";
		wait for Clk_period;
		Addr <=  "00110000101111";
		Trees_din <= x"03fd6504";
		wait for Clk_period;
		Addr <=  "00110000110000";
		Trees_din <= x"001930f5";
		wait for Clk_period;
		Addr <=  "00110000110001";
		Trees_din <= x"006330f5";
		wait for Clk_period;
		Addr <=  "00110000110010";
		Trees_din <= x"fff030f5";
		wait for Clk_period;
		Addr <=  "00110000110011";
		Trees_din <= x"0f01eb08";
		wait for Clk_period;
		Addr <=  "00110000110100";
		Trees_din <= x"09005104";
		wait for Clk_period;
		Addr <=  "00110000110101";
		Trees_din <= x"ff9830f5";
		wait for Clk_period;
		Addr <=  "00110000110110";
		Trees_din <= x"003430f5";
		wait for Clk_period;
		Addr <=  "00110000110111";
		Trees_din <= x"05fa7504";
		wait for Clk_period;
		Addr <=  "00110000111000";
		Trees_din <= x"004930f5";
		wait for Clk_period;
		Addr <=  "00110000111001";
		Trees_din <= x"ffdd30f5";
		wait for Clk_period;
		Addr <=  "00110000111010";
		Trees_din <= x"17002f04";
		wait for Clk_period;
		Addr <=  "00110000111011";
		Trees_din <= x"fffa30f5";
		wait for Clk_period;
		Addr <=  "00110000111100";
		Trees_din <= x"007a30f5";
		wait for Clk_period;
		Addr <=  "00110000111101";
		Trees_din <= x"000ceb3c";
		wait for Clk_period;
		Addr <=  "00110000111110";
		Trees_din <= x"08034328";
		wait for Clk_period;
		Addr <=  "00110000111111";
		Trees_din <= x"03f89814";
		wait for Clk_period;
		Addr <=  "00110001000000";
		Trees_din <= x"000b9b10";
		wait for Clk_period;
		Addr <=  "00110001000001";
		Trees_din <= x"0009b108";
		wait for Clk_period;
		Addr <=  "00110001000010";
		Trees_din <= x"14013504";
		wait for Clk_period;
		Addr <=  "00110001000011";
		Trees_din <= x"ffff31e1";
		wait for Clk_period;
		Addr <=  "00110001000100";
		Trees_din <= x"005631e1";
		wait for Clk_period;
		Addr <=  "00110001000101";
		Trees_din <= x"05fa0504";
		wait for Clk_period;
		Addr <=  "00110001000110";
		Trees_din <= x"001f31e1";
		wait for Clk_period;
		Addr <=  "00110001000111";
		Trees_din <= x"ffac31e1";
		wait for Clk_period;
		Addr <=  "00110001001000";
		Trees_din <= x"007a31e1";
		wait for Clk_period;
		Addr <=  "00110001001001";
		Trees_din <= x"01107310";
		wait for Clk_period;
		Addr <=  "00110001001010";
		Trees_din <= x"21000108";
		wait for Clk_period;
		Addr <=  "00110001001011";
		Trees_din <= x"07005e04";
		wait for Clk_period;
		Addr <=  "00110001001100";
		Trees_din <= x"000731e1";
		wait for Clk_period;
		Addr <=  "00110001001101";
		Trees_din <= x"ffb231e1";
		wait for Clk_period;
		Addr <=  "00110001001110";
		Trees_din <= x"05faba04";
		wait for Clk_period;
		Addr <=  "00110001001111";
		Trees_din <= x"006731e1";
		wait for Clk_period;
		Addr <=  "00110001010000";
		Trees_din <= x"000431e1";
		wait for Clk_period;
		Addr <=  "00110001010001";
		Trees_din <= x"ffa031e1";
		wait for Clk_period;
		Addr <=  "00110001010010";
		Trees_din <= x"0700540c";
		wait for Clk_period;
		Addr <=  "00110001010011";
		Trees_din <= x"1500ae08";
		wait for Clk_period;
		Addr <=  "00110001010100";
		Trees_din <= x"09005004";
		wait for Clk_period;
		Addr <=  "00110001010101";
		Trees_din <= x"ffe031e1";
		wait for Clk_period;
		Addr <=  "00110001010110";
		Trees_din <= x"000931e1";
		wait for Clk_period;
		Addr <=  "00110001010111";
		Trees_din <= x"005e31e1";
		wait for Clk_period;
		Addr <=  "00110001011000";
		Trees_din <= x"020abe04";
		wait for Clk_period;
		Addr <=  "00110001011001";
		Trees_din <= x"ff8d31e1";
		wait for Clk_period;
		Addr <=  "00110001011010";
		Trees_din <= x"fff831e1";
		wait for Clk_period;
		Addr <=  "00110001011011";
		Trees_din <= x"0803b638";
		wait for Clk_period;
		Addr <=  "00110001011100";
		Trees_din <= x"0d024f18";
		wait for Clk_period;
		Addr <=  "00110001011101";
		Trees_din <= x"0f03f610";
		wait for Clk_period;
		Addr <=  "00110001011110";
		Trees_din <= x"08020d08";
		wait for Clk_period;
		Addr <=  "00110001011111";
		Trees_din <= x"0afb1804";
		wait for Clk_period;
		Addr <=  "00110001100000";
		Trees_din <= x"ffe731e1";
		wait for Clk_period;
		Addr <=  "00110001100001";
		Trees_din <= x"ff8a31e1";
		wait for Clk_period;
		Addr <=  "00110001100010";
		Trees_din <= x"10028804";
		wait for Clk_period;
		Addr <=  "00110001100011";
		Trees_din <= x"ffbe31e1";
		wait for Clk_period;
		Addr <=  "00110001100100";
		Trees_din <= x"003a31e1";
		wait for Clk_period;
		Addr <=  "00110001100101";
		Trees_din <= x"06f48704";
		wait for Clk_period;
		Addr <=  "00110001100110";
		Trees_din <= x"006031e1";
		wait for Clk_period;
		Addr <=  "00110001100111";
		Trees_din <= x"fff331e1";
		wait for Clk_period;
		Addr <=  "00110001101000";
		Trees_din <= x"0d032e10";
		wait for Clk_period;
		Addr <=  "00110001101001";
		Trees_din <= x"06f49108";
		wait for Clk_period;
		Addr <=  "00110001101010";
		Trees_din <= x"12013b04";
		wait for Clk_period;
		Addr <=  "00110001101011";
		Trees_din <= x"ffaa31e1";
		wait for Clk_period;
		Addr <=  "00110001101100";
		Trees_din <= x"000d31e1";
		wait for Clk_period;
		Addr <=  "00110001101101";
		Trees_din <= x"0afb4704";
		wait for Clk_period;
		Addr <=  "00110001101110";
		Trees_din <= x"ffe731e1";
		wait for Clk_period;
		Addr <=  "00110001101111";
		Trees_din <= x"006931e1";
		wait for Clk_period;
		Addr <=  "00110001110000";
		Trees_din <= x"0af7f108";
		wait for Clk_period;
		Addr <=  "00110001110001";
		Trees_din <= x"0af7a504";
		wait for Clk_period;
		Addr <=  "00110001110010";
		Trees_din <= x"ffdb31e1";
		wait for Clk_period;
		Addr <=  "00110001110011";
		Trees_din <= x"007b31e1";
		wait for Clk_period;
		Addr <=  "00110001110100";
		Trees_din <= x"0f00c604";
		wait for Clk_period;
		Addr <=  "00110001110101";
		Trees_din <= x"ffe631e1";
		wait for Clk_period;
		Addr <=  "00110001110110";
		Trees_din <= x"ff8a31e1";
		wait for Clk_period;
		Addr <=  "00110001110111";
		Trees_din <= x"005631e1";
		wait for Clk_period;
		Addr <=  "00110001111000";
		Trees_din <= x"020baf58";
		wait for Clk_period;
		Addr <=  "00110001111001";
		Trees_din <= x"04f95824";
		wait for Clk_period;
		Addr <=  "00110001111010";
		Trees_din <= x"10f97c04";
		wait for Clk_period;
		Addr <=  "00110001111011";
		Trees_din <= x"ff9432f5";
		wait for Clk_period;
		Addr <=  "00110001111100";
		Trees_din <= x"0b028810";
		wait for Clk_period;
		Addr <=  "00110001111101";
		Trees_din <= x"0bfa8108";
		wait for Clk_period;
		Addr <=  "00110001111110";
		Trees_din <= x"1000f504";
		wait for Clk_period;
		Addr <=  "00110001111111";
		Trees_din <= x"005132f5";
		wait for Clk_period;
		Addr <=  "00110010000000";
		Trees_din <= x"ffcd32f5";
		wait for Clk_period;
		Addr <=  "00110010000001";
		Trees_din <= x"000d6304";
		wait for Clk_period;
		Addr <=  "00110010000010";
		Trees_din <= x"ffeb32f5";
		wait for Clk_period;
		Addr <=  "00110010000011";
		Trees_din <= x"ff9532f5";
		wait for Clk_period;
		Addr <=  "00110010000100";
		Trees_din <= x"1003ee08";
		wait for Clk_period;
		Addr <=  "00110010000101";
		Trees_din <= x"07005804";
		wait for Clk_period;
		Addr <=  "00110010000110";
		Trees_din <= x"001f32f5";
		wait for Clk_period;
		Addr <=  "00110010000111";
		Trees_din <= x"007432f5";
		wait for Clk_period;
		Addr <=  "00110010001000";
		Trees_din <= x"1f000004";
		wait for Clk_period;
		Addr <=  "00110010001001";
		Trees_din <= x"ffba32f5";
		wait for Clk_period;
		Addr <=  "00110010001010";
		Trees_din <= x"004e32f5";
		wait for Clk_period;
		Addr <=  "00110010001011";
		Trees_din <= x"0a03e220";
		wait for Clk_period;
		Addr <=  "00110010001100";
		Trees_din <= x"05fba710";
		wait for Clk_period;
		Addr <=  "00110010001101";
		Trees_din <= x"15009d08";
		wait for Clk_period;
		Addr <=  "00110010001110";
		Trees_din <= x"02ff5f04";
		wait for Clk_period;
		Addr <=  "00110010001111";
		Trees_din <= x"ffae32f5";
		wait for Clk_period;
		Addr <=  "00110010010000";
		Trees_din <= x"002a32f5";
		wait for Clk_period;
		Addr <=  "00110010010001";
		Trees_din <= x"04fe5b04";
		wait for Clk_period;
		Addr <=  "00110010010010";
		Trees_din <= x"001f32f5";
		wait for Clk_period;
		Addr <=  "00110010010011";
		Trees_din <= x"ffcd32f5";
		wait for Clk_period;
		Addr <=  "00110010010100";
		Trees_din <= x"0af7b408";
		wait for Clk_period;
		Addr <=  "00110010010101";
		Trees_din <= x"13fdbb04";
		wait for Clk_period;
		Addr <=  "00110010010110";
		Trees_din <= x"ff9232f5";
		wait for Clk_period;
		Addr <=  "00110010010111";
		Trees_din <= x"ffdb32f5";
		wait for Clk_period;
		Addr <=  "00110010011000";
		Trees_din <= x"02091304";
		wait for Clk_period;
		Addr <=  "00110010011001";
		Trees_din <= x"fff632f5";
		wait for Clk_period;
		Addr <=  "00110010011010";
		Trees_din <= x"003c32f5";
		wait for Clk_period;
		Addr <=  "00110010011011";
		Trees_din <= x"0d00da08";
		wait for Clk_period;
		Addr <=  "00110010011100";
		Trees_din <= x"19008f04";
		wait for Clk_period;
		Addr <=  "00110010011101";
		Trees_din <= x"ffbc32f5";
		wait for Clk_period;
		Addr <=  "00110010011110";
		Trees_din <= x"005432f5";
		wait for Clk_period;
		Addr <=  "00110010011111";
		Trees_din <= x"17000004";
		wait for Clk_period;
		Addr <=  "00110010100000";
		Trees_din <= x"001d32f5";
		wait for Clk_period;
		Addr <=  "00110010100001";
		Trees_din <= x"1b003104";
		wait for Clk_period;
		Addr <=  "00110010100010";
		Trees_din <= x"ffe632f5";
		wait for Clk_period;
		Addr <=  "00110010100011";
		Trees_din <= x"ff7e32f5";
		wait for Clk_period;
		Addr <=  "00110010100100";
		Trees_din <= x"1601120c";
		wait for Clk_period;
		Addr <=  "00110010100101";
		Trees_din <= x"13fd9808";
		wait for Clk_period;
		Addr <=  "00110010100110";
		Trees_din <= x"13f9d204";
		wait for Clk_period;
		Addr <=  "00110010100111";
		Trees_din <= x"004332f5";
		wait for Clk_period;
		Addr <=  "00110010101000";
		Trees_din <= x"ffbc32f5";
		wait for Clk_period;
		Addr <=  "00110010101001";
		Trees_din <= x"006c32f5";
		wait for Clk_period;
		Addr <=  "00110010101010";
		Trees_din <= x"17000d0c";
		wait for Clk_period;
		Addr <=  "00110010101011";
		Trees_din <= x"09005404";
		wait for Clk_period;
		Addr <=  "00110010101100";
		Trees_din <= x"001532f5";
		wait for Clk_period;
		Addr <=  "00110010101101";
		Trees_din <= x"04fb8704";
		wait for Clk_period;
		Addr <=  "00110010101110";
		Trees_din <= x"ff8f32f5";
		wait for Clk_period;
		Addr <=  "00110010101111";
		Trees_din <= x"ffee32f5";
		wait for Clk_period;
		Addr <=  "00110010110000";
		Trees_din <= x"1500990c";
		wait for Clk_period;
		Addr <=  "00110010110001";
		Trees_din <= x"14000d04";
		wait for Clk_period;
		Addr <=  "00110010110010";
		Trees_din <= x"ffd532f5";
		wait for Clk_period;
		Addr <=  "00110010110011";
		Trees_din <= x"11ff1104";
		wait for Clk_period;
		Addr <=  "00110010110100";
		Trees_din <= x"ffe832f5";
		wait for Clk_period;
		Addr <=  "00110010110101";
		Trees_din <= x"005d32f5";
		wait for Clk_period;
		Addr <=  "00110010110110";
		Trees_din <= x"1c002b08";
		wait for Clk_period;
		Addr <=  "00110010110111";
		Trees_din <= x"05fad804";
		wait for Clk_period;
		Addr <=  "00110010111000";
		Trees_din <= x"000632f5";
		wait for Clk_period;
		Addr <=  "00110010111001";
		Trees_din <= x"005d32f5";
		wait for Clk_period;
		Addr <=  "00110010111010";
		Trees_din <= x"13fe4804";
		wait for Clk_period;
		Addr <=  "00110010111011";
		Trees_din <= x"001d32f5";
		wait for Clk_period;
		Addr <=  "00110010111100";
		Trees_din <= x"ff9832f5";
		wait for Clk_period;
		Addr <=  "00110010111101";
		Trees_din <= x"1104aa58";
		wait for Clk_period;
		Addr <=  "00110010111110";
		Trees_din <= x"0c020b2c";
		wait for Clk_period;
		Addr <=  "00110010111111";
		Trees_din <= x"08028d1c";
		wait for Clk_period;
		Addr <=  "00110011000000";
		Trees_din <= x"0201230c";
		wait for Clk_period;
		Addr <=  "00110011000001";
		Trees_din <= x"08006404";
		wait for Clk_period;
		Addr <=  "00110011000010";
		Trees_din <= x"ff8b33b1";
		wait for Clk_period;
		Addr <=  "00110011000011";
		Trees_din <= x"0b04dc04";
		wait for Clk_period;
		Addr <=  "00110011000100";
		Trees_din <= x"ffda33b1";
		wait for Clk_period;
		Addr <=  "00110011000101";
		Trees_din <= x"003c33b1";
		wait for Clk_period;
		Addr <=  "00110011000110";
		Trees_din <= x"09005608";
		wait for Clk_period;
		Addr <=  "00110011000111";
		Trees_din <= x"0b028604";
		wait for Clk_period;
		Addr <=  "00110011001000";
		Trees_din <= x"002e33b1";
		wait for Clk_period;
		Addr <=  "00110011001001";
		Trees_din <= x"ffff33b1";
		wait for Clk_period;
		Addr <=  "00110011001010";
		Trees_din <= x"0c014c04";
		wait for Clk_period;
		Addr <=  "00110011001011";
		Trees_din <= x"000b33b1";
		wait for Clk_period;
		Addr <=  "00110011001100";
		Trees_din <= x"ffbc33b1";
		wait for Clk_period;
		Addr <=  "00110011001101";
		Trees_din <= x"0304d30c";
		wait for Clk_period;
		Addr <=  "00110011001110";
		Trees_din <= x"21000008";
		wait for Clk_period;
		Addr <=  "00110011001111";
		Trees_din <= x"1a00e304";
		wait for Clk_period;
		Addr <=  "00110011010000";
		Trees_din <= x"ff8a33b1";
		wait for Clk_period;
		Addr <=  "00110011010001";
		Trees_din <= x"ffe033b1";
		wait for Clk_period;
		Addr <=  "00110011010010";
		Trees_din <= x"002a33b1";
		wait for Clk_period;
		Addr <=  "00110011010011";
		Trees_din <= x"002a33b1";
		wait for Clk_period;
		Addr <=  "00110011010100";
		Trees_din <= x"09004c0c";
		wait for Clk_period;
		Addr <=  "00110011010101";
		Trees_din <= x"06f46e04";
		wait for Clk_period;
		Addr <=  "00110011010110";
		Trees_din <= x"000b33b1";
		wait for Clk_period;
		Addr <=  "00110011010111";
		Trees_din <= x"0800e704";
		wait for Clk_period;
		Addr <=  "00110011011000";
		Trees_din <= x"ffe433b1";
		wait for Clk_period;
		Addr <=  "00110011011001";
		Trees_din <= x"ff8d33b1";
		wait for Clk_period;
		Addr <=  "00110011011010";
		Trees_din <= x"0c02c510";
		wait for Clk_period;
		Addr <=  "00110011011011";
		Trees_din <= x"07005908";
		wait for Clk_period;
		Addr <=  "00110011011100";
		Trees_din <= x"0d036804";
		wait for Clk_period;
		Addr <=  "00110011011101";
		Trees_din <= x"002033b1";
		wait for Clk_period;
		Addr <=  "00110011011110";
		Trees_din <= x"ffc133b1";
		wait for Clk_period;
		Addr <=  "00110011011111";
		Trees_din <= x"0203a104";
		wait for Clk_period;
		Addr <=  "00110011100000";
		Trees_din <= x"ffff33b1";
		wait for Clk_period;
		Addr <=  "00110011100001";
		Trees_din <= x"006f33b1";
		wait for Clk_period;
		Addr <=  "00110011100010";
		Trees_din <= x"04fff308";
		wait for Clk_period;
		Addr <=  "00110011100011";
		Trees_din <= x"0f00c604";
		wait for Clk_period;
		Addr <=  "00110011100100";
		Trees_din <= x"001a33b1";
		wait for Clk_period;
		Addr <=  "00110011100101";
		Trees_din <= x"ffc333b1";
		wait for Clk_period;
		Addr <=  "00110011100110";
		Trees_din <= x"00021604";
		wait for Clk_period;
		Addr <=  "00110011100111";
		Trees_din <= x"fffa33b1";
		wait for Clk_period;
		Addr <=  "00110011101000";
		Trees_din <= x"004a33b1";
		wait for Clk_period;
		Addr <=  "00110011101001";
		Trees_din <= x"09005504";
		wait for Clk_period;
		Addr <=  "00110011101010";
		Trees_din <= x"fff933b1";
		wait for Clk_period;
		Addr <=  "00110011101011";
		Trees_din <= x"ffab33b1";
		wait for Clk_period;
		Addr <=  "00110011101100";
		Trees_din <= x"020b6158";
		wait for Clk_period;
		Addr <=  "00110011101101";
		Trees_din <= x"04fa4d2c";
		wait for Clk_period;
		Addr <=  "00110011101110";
		Trees_din <= x"0bfa8114";
		wait for Clk_period;
		Addr <=  "00110011101111";
		Trees_din <= x"0bf9c710";
		wait for Clk_period;
		Addr <=  "00110011110000";
		Trees_din <= x"14011708";
		wait for Clk_period;
		Addr <=  "00110011110001";
		Trees_din <= x"03f70404";
		wait for Clk_period;
		Addr <=  "00110011110010";
		Trees_din <= x"ffea34b5";
		wait for Clk_period;
		Addr <=  "00110011110011";
		Trees_din <= x"004434b5";
		wait for Clk_period;
		Addr <=  "00110011110100";
		Trees_din <= x"12021004";
		wait for Clk_period;
		Addr <=  "00110011110101";
		Trees_din <= x"ffaa34b5";
		wait for Clk_period;
		Addr <=  "00110011110110";
		Trees_din <= x"fffb34b5";
		wait for Clk_period;
		Addr <=  "00110011110111";
		Trees_din <= x"004b34b5";
		wait for Clk_period;
		Addr <=  "00110011111000";
		Trees_din <= x"04f4e308";
		wait for Clk_period;
		Addr <=  "00110011111001";
		Trees_din <= x"04f47104";
		wait for Clk_period;
		Addr <=  "00110011111010";
		Trees_din <= x"ffe034b5";
		wait for Clk_period;
		Addr <=  "00110011111011";
		Trees_din <= x"005934b5";
		wait for Clk_period;
		Addr <=  "00110011111100";
		Trees_din <= x"18003908";
		wait for Clk_period;
		Addr <=  "00110011111101";
		Trees_din <= x"03f89804";
		wait for Clk_period;
		Addr <=  "00110011111110";
		Trees_din <= x"004234b5";
		wait for Clk_period;
		Addr <=  "00110011111111";
		Trees_din <= x"ffc934b5";
		wait for Clk_period;
		Addr <=  "00110100000000";
		Trees_din <= x"18004804";
		wait for Clk_period;
		Addr <=  "00110100000001";
		Trees_din <= x"ff9334b5";
		wait for Clk_period;
		Addr <=  "00110100000010";
		Trees_din <= x"fff034b5";
		wait for Clk_period;
		Addr <=  "00110100000011";
		Trees_din <= x"06f8921c";
		wait for Clk_period;
		Addr <=  "00110100000100";
		Trees_din <= x"19009e10";
		wait for Clk_period;
		Addr <=  "00110100000101";
		Trees_din <= x"19009b08";
		wait for Clk_period;
		Addr <=  "00110100000110";
		Trees_din <= x"0c02dd04";
		wait for Clk_period;
		Addr <=  "00110100000111";
		Trees_din <= x"000a34b5";
		wait for Clk_period;
		Addr <=  "00110100001000";
		Trees_din <= x"ffd834b5";
		wait for Clk_period;
		Addr <=  "00110100001001";
		Trees_din <= x"06f39904";
		wait for Clk_period;
		Addr <=  "00110100001010";
		Trees_din <= x"ffe634b5";
		wait for Clk_period;
		Addr <=  "00110100001011";
		Trees_din <= x"005534b5";
		wait for Clk_period;
		Addr <=  "00110100001100";
		Trees_din <= x"15009304";
		wait for Clk_period;
		Addr <=  "00110100001101";
		Trees_din <= x"ff9434b5";
		wait for Clk_period;
		Addr <=  "00110100001110";
		Trees_din <= x"02079804";
		wait for Clk_period;
		Addr <=  "00110100001111";
		Trees_din <= x"ffdf34b5";
		wait for Clk_period;
		Addr <=  "00110100010000";
		Trees_din <= x"002534b5";
		wait for Clk_period;
		Addr <=  "00110100010001";
		Trees_din <= x"11fecd04";
		wait for Clk_period;
		Addr <=  "00110100010010";
		Trees_din <= x"ffae34b5";
		wait for Clk_period;
		Addr <=  "00110100010011";
		Trees_din <= x"0f001f04";
		wait for Clk_period;
		Addr <=  "00110100010100";
		Trees_din <= x"ffcb34b5";
		wait for Clk_period;
		Addr <=  "00110100010101";
		Trees_din <= x"1e005904";
		wait for Clk_period;
		Addr <=  "00110100010110";
		Trees_din <= x"fff534b5";
		wait for Clk_period;
		Addr <=  "00110100010111";
		Trees_din <= x"005934b5";
		wait for Clk_period;
		Addr <=  "00110100011000";
		Trees_din <= x"0700530c";
		wait for Clk_period;
		Addr <=  "00110100011001";
		Trees_din <= x"06f3df08";
		wait for Clk_period;
		Addr <=  "00110100011010";
		Trees_din <= x"17002904";
		wait for Clk_period;
		Addr <=  "00110100011011";
		Trees_din <= x"ffd434b5";
		wait for Clk_period;
		Addr <=  "00110100011100";
		Trees_din <= x"002e34b5";
		wait for Clk_period;
		Addr <=  "00110100011101";
		Trees_din <= x"006334b5";
		wait for Clk_period;
		Addr <=  "00110100011110";
		Trees_din <= x"1601120c";
		wait for Clk_period;
		Addr <=  "00110100011111";
		Trees_din <= x"13fd9808";
		wait for Clk_period;
		Addr <=  "00110100100000";
		Trees_din <= x"13f9e204";
		wait for Clk_period;
		Addr <=  "00110100100001";
		Trees_din <= x"002334b5";
		wait for Clk_period;
		Addr <=  "00110100100010";
		Trees_din <= x"ffcc34b5";
		wait for Clk_period;
		Addr <=  "00110100100011";
		Trees_din <= x"006834b5";
		wait for Clk_period;
		Addr <=  "00110100100100";
		Trees_din <= x"1c00420c";
		wait for Clk_period;
		Addr <=  "00110100100101";
		Trees_din <= x"0003e504";
		wait for Clk_period;
		Addr <=  "00110100100110";
		Trees_din <= x"004e34b5";
		wait for Clk_period;
		Addr <=  "00110100100111";
		Trees_din <= x"05fc8504";
		wait for Clk_period;
		Addr <=  "00110100101000";
		Trees_din <= x"ffb834b5";
		wait for Clk_period;
		Addr <=  "00110100101001";
		Trees_din <= x"000034b5";
		wait for Clk_period;
		Addr <=  "00110100101010";
		Trees_din <= x"09005404";
		wait for Clk_period;
		Addr <=  "00110100101011";
		Trees_din <= x"fff934b5";
		wait for Clk_period;
		Addr <=  "00110100101100";
		Trees_din <= x"005c34b5";
		wait for Clk_period;
		Addr <=  "00110100101101";
		Trees_din <= x"020c6044";
		wait for Clk_period;
		Addr <=  "00110100101110";
		Trees_din <= x"03f44a04";
		wait for Clk_period;
		Addr <=  "00110100101111";
		Trees_din <= x"ffb53589";
		wait for Clk_period;
		Addr <=  "00110100110000";
		Trees_din <= x"0f000420";
		wait for Clk_period;
		Addr <=  "00110100110001";
		Trees_din <= x"1200da10";
		wait for Clk_period;
		Addr <=  "00110100110010";
		Trees_din <= x"12ff0f08";
		wait for Clk_period;
		Addr <=  "00110100110011";
		Trees_din <= x"10050804";
		wait for Clk_period;
		Addr <=  "00110100110100";
		Trees_din <= x"ffd13589";
		wait for Clk_period;
		Addr <=  "00110100110101";
		Trees_din <= x"002f3589";
		wait for Clk_period;
		Addr <=  "00110100110110";
		Trees_din <= x"0c012004";
		wait for Clk_period;
		Addr <=  "00110100110111";
		Trees_din <= x"00783589";
		wait for Clk_period;
		Addr <=  "00110100111000";
		Trees_din <= x"000a3589";
		wait for Clk_period;
		Addr <=  "00110100111001";
		Trees_din <= x"14010408";
		wait for Clk_period;
		Addr <=  "00110100111010";
		Trees_din <= x"1703ac04";
		wait for Clk_period;
		Addr <=  "00110100111011";
		Trees_din <= x"ffab3589";
		wait for Clk_period;
		Addr <=  "00110100111100";
		Trees_din <= x"00133589";
		wait for Clk_period;
		Addr <=  "00110100111101";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00110100111110";
		Trees_din <= x"004f3589";
		wait for Clk_period;
		Addr <=  "00110100111111";
		Trees_din <= x"ffc23589";
		wait for Clk_period;
		Addr <=  "00110101000000";
		Trees_din <= x"17012b10";
		wait for Clk_period;
		Addr <=  "00110101000001";
		Trees_din <= x"1700eb08";
		wait for Clk_period;
		Addr <=  "00110101000010";
		Trees_din <= x"1b003004";
		wait for Clk_period;
		Addr <=  "00110101000011";
		Trees_din <= x"ffcd3589";
		wait for Clk_period;
		Addr <=  "00110101000100";
		Trees_din <= x"00073589";
		wait for Clk_period;
		Addr <=  "00110101000101";
		Trees_din <= x"1400d904";
		wait for Clk_period;
		Addr <=  "00110101000110";
		Trees_din <= x"ffee3589";
		wait for Clk_period;
		Addr <=  "00110101000111";
		Trees_din <= x"005d3589";
		wait for Clk_period;
		Addr <=  "00110101001000";
		Trees_din <= x"0afccc08";
		wait for Clk_period;
		Addr <=  "00110101001001";
		Trees_din <= x"1200ae04";
		wait for Clk_period;
		Addr <=  "00110101001010";
		Trees_din <= x"ffa73589";
		wait for Clk_period;
		Addr <=  "00110101001011";
		Trees_din <= x"00123589";
		wait for Clk_period;
		Addr <=  "00110101001100";
		Trees_din <= x"12fe4404";
		wait for Clk_period;
		Addr <=  "00110101001101";
		Trees_din <= x"00133589";
		wait for Clk_period;
		Addr <=  "00110101001110";
		Trees_din <= x"ffb43589";
		wait for Clk_period;
		Addr <=  "00110101001111";
		Trees_din <= x"00037704";
		wait for Clk_period;
		Addr <=  "00110101010000";
		Trees_din <= x"00643589";
		wait for Clk_period;
		Addr <=  "00110101010001";
		Trees_din <= x"0f000b08";
		wait for Clk_period;
		Addr <=  "00110101010010";
		Trees_din <= x"05fb8404";
		wait for Clk_period;
		Addr <=  "00110101010011";
		Trees_din <= x"ffaf3589";
		wait for Clk_period;
		Addr <=  "00110101010100";
		Trees_din <= x"00223589";
		wait for Clk_period;
		Addr <=  "00110101010101";
		Trees_din <= x"17000d10";
		wait for Clk_period;
		Addr <=  "00110101010110";
		Trees_din <= x"16011208";
		wait for Clk_period;
		Addr <=  "00110101010111";
		Trees_din <= x"13fd9804";
		wait for Clk_period;
		Addr <=  "00110101011000";
		Trees_din <= x"ffe93589";
		wait for Clk_period;
		Addr <=  "00110101011001";
		Trees_din <= x"00513589";
		wait for Clk_period;
		Addr <=  "00110101011010";
		Trees_din <= x"09005604";
		wait for Clk_period;
		Addr <=  "00110101011011";
		Trees_din <= x"ffe23589";
		wait for Clk_period;
		Addr <=  "00110101011100";
		Trees_din <= x"ff9e3589";
		wait for Clk_period;
		Addr <=  "00110101011101";
		Trees_din <= x"12fef604";
		wait for Clk_period;
		Addr <=  "00110101011110";
		Trees_din <= x"ffe13589";
		wait for Clk_period;
		Addr <=  "00110101011111";
		Trees_din <= x"02112404";
		wait for Clk_period;
		Addr <=  "00110101100000";
		Trees_din <= x"00583589";
		wait for Clk_period;
		Addr <=  "00110101100001";
		Trees_din <= x"fff53589";
		wait for Clk_period;
		Addr <=  "00110101100010";
		Trees_din <= x"02047558";
		wait for Clk_period;
		Addr <=  "00110101100011";
		Trees_din <= x"0402ed30";
		wait for Clk_period;
		Addr <=  "00110101100100";
		Trees_din <= x"07005518";
		wait for Clk_period;
		Addr <=  "00110101100101";
		Trees_din <= x"1202810c";
		wait for Clk_period;
		Addr <=  "00110101100110";
		Trees_din <= x"08017008";
		wait for Clk_period;
		Addr <=  "00110101100111";
		Trees_din <= x"08007604";
		wait for Clk_period;
		Addr <=  "00110101101000";
		Trees_din <= x"ffb436c5";
		wait for Clk_period;
		Addr <=  "00110101101001";
		Trees_din <= x"003f36c5";
		wait for Clk_period;
		Addr <=  "00110101101010";
		Trees_din <= x"ff9636c5";
		wait for Clk_period;
		Addr <=  "00110101101011";
		Trees_din <= x"0801cf04";
		wait for Clk_period;
		Addr <=  "00110101101100";
		Trees_din <= x"ffdc36c5";
		wait for Clk_period;
		Addr <=  "00110101101101";
		Trees_din <= x"0d015a04";
		wait for Clk_period;
		Addr <=  "00110101101110";
		Trees_din <= x"001636c5";
		wait for Clk_period;
		Addr <=  "00110101101111";
		Trees_din <= x"007636c5";
		wait for Clk_period;
		Addr <=  "00110101110000";
		Trees_din <= x"05f89e08";
		wait for Clk_period;
		Addr <=  "00110101110001";
		Trees_din <= x"09005904";
		wait for Clk_period;
		Addr <=  "00110101110010";
		Trees_din <= x"fff036c5";
		wait for Clk_period;
		Addr <=  "00110101110011";
		Trees_din <= x"005b36c5";
		wait for Clk_period;
		Addr <=  "00110101110100";
		Trees_din <= x"06f84408";
		wait for Clk_period;
		Addr <=  "00110101110101";
		Trees_din <= x"13f90f04";
		wait for Clk_period;
		Addr <=  "00110101110110";
		Trees_din <= x"ffe836c5";
		wait for Clk_period;
		Addr <=  "00110101110111";
		Trees_din <= x"ff8336c5";
		wait for Clk_period;
		Addr <=  "00110101111000";
		Trees_din <= x"0afb2b04";
		wait for Clk_period;
		Addr <=  "00110101111001";
		Trees_din <= x"002c36c5";
		wait for Clk_period;
		Addr <=  "00110101111010";
		Trees_din <= x"ffbf36c5";
		wait for Clk_period;
		Addr <=  "00110101111011";
		Trees_din <= x"0406be18";
		wait for Clk_period;
		Addr <=  "00110101111100";
		Trees_din <= x"1102840c";
		wait for Clk_period;
		Addr <=  "00110101111101";
		Trees_din <= x"01087508";
		wait for Clk_period;
		Addr <=  "00110101111110";
		Trees_din <= x"0f009f04";
		wait for Clk_period;
		Addr <=  "00110101111111";
		Trees_din <= x"000c36c5";
		wait for Clk_period;
		Addr <=  "00110110000000";
		Trees_din <= x"005b36c5";
		wait for Clk_period;
		Addr <=  "00110110000001";
		Trees_din <= x"ffdf36c5";
		wait for Clk_period;
		Addr <=  "00110110000010";
		Trees_din <= x"07005908";
		wait for Clk_period;
		Addr <=  "00110110000011";
		Trees_din <= x"02013704";
		wait for Clk_period;
		Addr <=  "00110110000100";
		Trees_din <= x"ffa236c5";
		wait for Clk_period;
		Addr <=  "00110110000101";
		Trees_din <= x"fff536c5";
		wait for Clk_period;
		Addr <=  "00110110000110";
		Trees_din <= x"003836c5";
		wait for Clk_period;
		Addr <=  "00110110000111";
		Trees_din <= x"1a009e04";
		wait for Clk_period;
		Addr <=  "00110110001000";
		Trees_din <= x"002336c5";
		wait for Clk_period;
		Addr <=  "00110110001001";
		Trees_din <= x"17001704";
		wait for Clk_period;
		Addr <=  "00110110001010";
		Trees_din <= x"ff8f36c5";
		wait for Clk_period;
		Addr <=  "00110110001011";
		Trees_din <= x"06f44e04";
		wait for Clk_period;
		Addr <=  "00110110001100";
		Trees_din <= x"002a36c5";
		wait for Clk_period;
		Addr <=  "00110110001101";
		Trees_din <= x"ffc536c5";
		wait for Clk_period;
		Addr <=  "00110110001110";
		Trees_din <= x"10f9731c";
		wait for Clk_period;
		Addr <=  "00110110001111";
		Trees_din <= x"04fbba0c";
		wait for Clk_period;
		Addr <=  "00110110010000";
		Trees_din <= x"01052804";
		wait for Clk_period;
		Addr <=  "00110110010001";
		Trees_din <= x"003a36c5";
		wait for Clk_period;
		Addr <=  "00110110010010";
		Trees_din <= x"15009c04";
		wait for Clk_period;
		Addr <=  "00110110010011";
		Trees_din <= x"ff9736c5";
		wait for Clk_period;
		Addr <=  "00110110010100";
		Trees_din <= x"fff236c5";
		wait for Clk_period;
		Addr <=  "00110110010101";
		Trees_din <= x"06f3d608";
		wait for Clk_period;
		Addr <=  "00110110010110";
		Trees_din <= x"05fa9f04";
		wait for Clk_period;
		Addr <=  "00110110010111";
		Trees_din <= x"ffd536c5";
		wait for Clk_period;
		Addr <=  "00110110011000";
		Trees_din <= x"003236c5";
		wait for Clk_period;
		Addr <=  "00110110011001";
		Trees_din <= x"0d01c804";
		wait for Clk_period;
		Addr <=  "00110110011010";
		Trees_din <= x"fff336c5";
		wait for Clk_period;
		Addr <=  "00110110011011";
		Trees_din <= x"009736c5";
		wait for Clk_period;
		Addr <=  "00110110011100";
		Trees_din <= x"04f68010";
		wait for Clk_period;
		Addr <=  "00110110011101";
		Trees_din <= x"0014ad0c";
		wait for Clk_period;
		Addr <=  "00110110011110";
		Trees_din <= x"1004ba08";
		wait for Clk_period;
		Addr <=  "00110110011111";
		Trees_din <= x"18004704";
		wait for Clk_period;
		Addr <=  "00110110100000";
		Trees_din <= x"007236c5";
		wait for Clk_period;
		Addr <=  "00110110100001";
		Trees_din <= x"001536c5";
		wait for Clk_period;
		Addr <=  "00110110100010";
		Trees_din <= x"000136c5";
		wait for Clk_period;
		Addr <=  "00110110100011";
		Trees_din <= x"ffc936c5";
		wait for Clk_period;
		Addr <=  "00110110100100";
		Trees_din <= x"0c006e0c";
		wait for Clk_period;
		Addr <=  "00110110100101";
		Trees_din <= x"0f03fb08";
		wait for Clk_period;
		Addr <=  "00110110100110";
		Trees_din <= x"01038904";
		wait for Clk_period;
		Addr <=  "00110110100111";
		Trees_din <= x"fff736c5";
		wait for Clk_period;
		Addr <=  "00110110101000";
		Trees_din <= x"005836c5";
		wait for Clk_period;
		Addr <=  "00110110101001";
		Trees_din <= x"ffc536c5";
		wait for Clk_period;
		Addr <=  "00110110101010";
		Trees_din <= x"0c00ad08";
		wait for Clk_period;
		Addr <=  "00110110101011";
		Trees_din <= x"06f4d304";
		wait for Clk_period;
		Addr <=  "00110110101100";
		Trees_din <= x"ff9d36c5";
		wait for Clk_period;
		Addr <=  "00110110101101";
		Trees_din <= x"000e36c5";
		wait for Clk_period;
		Addr <=  "00110110101110";
		Trees_din <= x"0d00d104";
		wait for Clk_period;
		Addr <=  "00110110101111";
		Trees_din <= x"002336c5";
		wait for Clk_period;
		Addr <=  "00110110110000";
		Trees_din <= x"fff436c5";
		wait for Clk_period;
		Addr <=  "00110110110001";
		Trees_din <= x"02083234";
		wait for Clk_period;
		Addr <=  "00110110110010";
		Trees_din <= x"0c03d72c";
		wait for Clk_period;
		Addr <=  "00110110110011";
		Trees_din <= x"07005314";
		wait for Clk_period;
		Addr <=  "00110110110100";
		Trees_din <= x"16001204";
		wait for Clk_period;
		Addr <=  "00110110110101";
		Trees_din <= x"005e37b9";
		wait for Clk_period;
		Addr <=  "00110110110110";
		Trees_din <= x"1c002708";
		wait for Clk_period;
		Addr <=  "00110110110111";
		Trees_din <= x"04012004";
		wait for Clk_period;
		Addr <=  "00110110111000";
		Trees_din <= x"ffcf37b9";
		wait for Clk_period;
		Addr <=  "00110110111001";
		Trees_din <= x"004337b9";
		wait for Clk_period;
		Addr <=  "00110110111010";
		Trees_din <= x"0c02dd04";
		wait for Clk_period;
		Addr <=  "00110110111011";
		Trees_din <= x"ff9737b9";
		wait for Clk_period;
		Addr <=  "00110110111100";
		Trees_din <= x"001137b9";
		wait for Clk_period;
		Addr <=  "00110110111101";
		Trees_din <= x"0f03f710";
		wait for Clk_period;
		Addr <=  "00110110111110";
		Trees_din <= x"0d000e08";
		wait for Clk_period;
		Addr <=  "00110110111111";
		Trees_din <= x"0c00e304";
		wait for Clk_period;
		Addr <=  "00110111000000";
		Trees_din <= x"006537b9";
		wait for Clk_period;
		Addr <=  "00110111000001";
		Trees_din <= x"fff337b9";
		wait for Clk_period;
		Addr <=  "00110111000010";
		Trees_din <= x"07005304";
		wait for Clk_period;
		Addr <=  "00110111000011";
		Trees_din <= x"005937b9";
		wait for Clk_period;
		Addr <=  "00110111000100";
		Trees_din <= x"fffe37b9";
		wait for Clk_period;
		Addr <=  "00110111000101";
		Trees_din <= x"01020f04";
		wait for Clk_period;
		Addr <=  "00110111000110";
		Trees_din <= x"000137b9";
		wait for Clk_period;
		Addr <=  "00110111000111";
		Trees_din <= x"ff8f37b9";
		wait for Clk_period;
		Addr <=  "00110111001000";
		Trees_din <= x"01049604";
		wait for Clk_period;
		Addr <=  "00110111001001";
		Trees_din <= x"fff637b9";
		wait for Clk_period;
		Addr <=  "00110111001010";
		Trees_din <= x"ffaa37b9";
		wait for Clk_period;
		Addr <=  "00110111001011";
		Trees_din <= x"1b004430";
		wait for Clk_period;
		Addr <=  "00110111001100";
		Trees_din <= x"0b028714";
		wait for Clk_period;
		Addr <=  "00110111001101";
		Trees_din <= x"10f9f904";
		wait for Clk_period;
		Addr <=  "00110111001110";
		Trees_din <= x"004e37b9";
		wait for Clk_period;
		Addr <=  "00110111001111";
		Trees_din <= x"0a017108";
		wait for Clk_period;
		Addr <=  "00110111010000";
		Trees_din <= x"0c01a204";
		wait for Clk_period;
		Addr <=  "00110111010001";
		Trees_din <= x"003037b9";
		wait for Clk_period;
		Addr <=  "00110111010010";
		Trees_din <= x"ffee37b9";
		wait for Clk_period;
		Addr <=  "00110111010011";
		Trees_din <= x"0f02fb04";
		wait for Clk_period;
		Addr <=  "00110111010100";
		Trees_din <= x"ffbf37b9";
		wait for Clk_period;
		Addr <=  "00110111010101";
		Trees_din <= x"001737b9";
		wait for Clk_period;
		Addr <=  "00110111010110";
		Trees_din <= x"04faa910";
		wait for Clk_period;
		Addr <=  "00110111010111";
		Trees_din <= x"0c026808";
		wait for Clk_period;
		Addr <=  "00110111011000";
		Trees_din <= x"09005904";
		wait for Clk_period;
		Addr <=  "00110111011001";
		Trees_din <= x"ffc237b9";
		wait for Clk_period;
		Addr <=  "00110111011010";
		Trees_din <= x"002d37b9";
		wait for Clk_period;
		Addr <=  "00110111011011";
		Trees_din <= x"0d031e04";
		wait for Clk_period;
		Addr <=  "00110111011100";
		Trees_din <= x"005a37b9";
		wait for Clk_period;
		Addr <=  "00110111011101";
		Trees_din <= x"000037b9";
		wait for Clk_period;
		Addr <=  "00110111011110";
		Trees_din <= x"1603f408";
		wait for Clk_period;
		Addr <=  "00110111011111";
		Trees_din <= x"0e01da04";
		wait for Clk_period;
		Addr <=  "00110111100000";
		Trees_din <= x"007037b9";
		wait for Clk_period;
		Addr <=  "00110111100001";
		Trees_din <= x"001337b9";
		wait for Clk_period;
		Addr <=  "00110111100010";
		Trees_din <= x"fffe37b9";
		wait for Clk_period;
		Addr <=  "00110111100011";
		Trees_din <= x"0a027610";
		wait for Clk_period;
		Addr <=  "00110111100100";
		Trees_din <= x"03f5fd04";
		wait for Clk_period;
		Addr <=  "00110111100101";
		Trees_din <= x"004537b9";
		wait for Clk_period;
		Addr <=  "00110111100110";
		Trees_din <= x"000f0708";
		wait for Clk_period;
		Addr <=  "00110111100111";
		Trees_din <= x"11023204";
		wait for Clk_period;
		Addr <=  "00110111101000";
		Trees_din <= x"ffdf37b9";
		wait for Clk_period;
		Addr <=  "00110111101001";
		Trees_din <= x"004737b9";
		wait for Clk_period;
		Addr <=  "00110111101010";
		Trees_din <= x"ffa837b9";
		wait for Clk_period;
		Addr <=  "00110111101011";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00110111101100";
		Trees_din <= x"ff9137b9";
		wait for Clk_period;
		Addr <=  "00110111101101";
		Trees_din <= x"fff237b9";
		wait for Clk_period;
		Addr <=  "00110111101110";
		Trees_din <= x"02047538";
		wait for Clk_period;
		Addr <=  "00110111101111";
		Trees_din <= x"16006510";
		wait for Clk_period;
		Addr <=  "00110111110000";
		Trees_din <= x"2100000c";
		wait for Clk_period;
		Addr <=  "00110111110001";
		Trees_din <= x"05fdec08";
		wait for Clk_period;
		Addr <=  "00110111110010";
		Trees_din <= x"19008204";
		wait for Clk_period;
		Addr <=  "00110111110011";
		Trees_din <= x"ffea38b5";
		wait for Clk_period;
		Addr <=  "00110111110100";
		Trees_din <= x"ff8938b5";
		wait for Clk_period;
		Addr <=  "00110111110101";
		Trees_din <= x"000738b5";
		wait for Clk_period;
		Addr <=  "00110111110110";
		Trees_din <= x"002338b5";
		wait for Clk_period;
		Addr <=  "00110111110111";
		Trees_din <= x"0a033220";
		wait for Clk_period;
		Addr <=  "00110111111000";
		Trees_din <= x"0d033710";
		wait for Clk_period;
		Addr <=  "00110111111001";
		Trees_din <= x"0d02e908";
		wait for Clk_period;
		Addr <=  "00110111111010";
		Trees_din <= x"0d02a704";
		wait for Clk_period;
		Addr <=  "00110111111011";
		Trees_din <= x"000c38b5";
		wait for Clk_period;
		Addr <=  "00110111111100";
		Trees_din <= x"ffad38b5";
		wait for Clk_period;
		Addr <=  "00110111111101";
		Trees_din <= x"05fd4e04";
		wait for Clk_period;
		Addr <=  "00110111111110";
		Trees_din <= x"005f38b5";
		wait for Clk_period;
		Addr <=  "00110111111111";
		Trees_din <= x"fff038b5";
		wait for Clk_period;
		Addr <=  "00111000000000";
		Trees_din <= x"1700f108";
		wait for Clk_period;
		Addr <=  "00111000000001";
		Trees_din <= x"08002d04";
		wait for Clk_period;
		Addr <=  "00111000000010";
		Trees_din <= x"000338b5";
		wait for Clk_period;
		Addr <=  "00111000000011";
		Trees_din <= x"ff8f38b5";
		wait for Clk_period;
		Addr <=  "00111000000100";
		Trees_din <= x"1b003e04";
		wait for Clk_period;
		Addr <=  "00111000000101";
		Trees_din <= x"ffe038b5";
		wait for Clk_period;
		Addr <=  "00111000000110";
		Trees_din <= x"004538b5";
		wait for Clk_period;
		Addr <=  "00111000000111";
		Trees_din <= x"0d014404";
		wait for Clk_period;
		Addr <=  "00111000001000";
		Trees_din <= x"fff738b5";
		wait for Clk_period;
		Addr <=  "00111000001001";
		Trees_din <= x"ff9b38b5";
		wait for Clk_period;
		Addr <=  "00111000001010";
		Trees_din <= x"00fe7b0c";
		wait for Clk_period;
		Addr <=  "00111000001011";
		Trees_din <= x"12ff0204";
		wait for Clk_period;
		Addr <=  "00111000001100";
		Trees_din <= x"fff238b5";
		wait for Clk_period;
		Addr <=  "00111000001101";
		Trees_din <= x"19008c04";
		wait for Clk_period;
		Addr <=  "00111000001110";
		Trees_din <= x"000638b5";
		wait for Clk_period;
		Addr <=  "00111000001111";
		Trees_din <= x"005838b5";
		wait for Clk_period;
		Addr <=  "00111000010000";
		Trees_din <= x"0bf9f61c";
		wait for Clk_period;
		Addr <=  "00111000010001";
		Trees_din <= x"1603db10";
		wait for Clk_period;
		Addr <=  "00111000010010";
		Trees_din <= x"08023808";
		wait for Clk_period;
		Addr <=  "00111000010011";
		Trees_din <= x"08005a04";
		wait for Clk_period;
		Addr <=  "00111000010100";
		Trees_din <= x"001138b5";
		wait for Clk_period;
		Addr <=  "00111000010101";
		Trees_din <= x"ffaa38b5";
		wait for Clk_period;
		Addr <=  "00111000010110";
		Trees_din <= x"07005604";
		wait for Clk_period;
		Addr <=  "00111000010111";
		Trees_din <= x"fff038b5";
		wait for Clk_period;
		Addr <=  "00111000011000";
		Trees_din <= x"004a38b5";
		wait for Clk_period;
		Addr <=  "00111000011001";
		Trees_din <= x"06f26204";
		wait for Clk_period;
		Addr <=  "00111000011010";
		Trees_din <= x"ffd938b5";
		wait for Clk_period;
		Addr <=  "00111000011011";
		Trees_din <= x"03f9a004";
		wait for Clk_period;
		Addr <=  "00111000011100";
		Trees_din <= x"002138b5";
		wait for Clk_period;
		Addr <=  "00111000011101";
		Trees_din <= x"006938b5";
		wait for Clk_period;
		Addr <=  "00111000011110";
		Trees_din <= x"0bfac510";
		wait for Clk_period;
		Addr <=  "00111000011111";
		Trees_din <= x"06f51308";
		wait for Clk_period;
		Addr <=  "00111000100000";
		Trees_din <= x"00097404";
		wait for Clk_period;
		Addr <=  "00111000100001";
		Trees_din <= x"002c38b5";
		wait for Clk_period;
		Addr <=  "00111000100010";
		Trees_din <= x"ffdf38b5";
		wait for Clk_period;
		Addr <=  "00111000100011";
		Trees_din <= x"02063404";
		wait for Clk_period;
		Addr <=  "00111000100100";
		Trees_din <= x"000938b5";
		wait for Clk_period;
		Addr <=  "00111000100101";
		Trees_din <= x"007338b5";
		wait for Clk_period;
		Addr <=  "00111000100110";
		Trees_din <= x"01029908";
		wait for Clk_period;
		Addr <=  "00111000100111";
		Trees_din <= x"14012704";
		wait for Clk_period;
		Addr <=  "00111000101000";
		Trees_din <= x"ffe838b5";
		wait for Clk_period;
		Addr <=  "00111000101001";
		Trees_din <= x"003d38b5";
		wait for Clk_period;
		Addr <=  "00111000101010";
		Trees_din <= x"05fc1804";
		wait for Clk_period;
		Addr <=  "00111000101011";
		Trees_din <= x"000638b5";
		wait for Clk_period;
		Addr <=  "00111000101100";
		Trees_din <= x"ffd038b5";
		wait for Clk_period;
		Addr <=  "00111000101101";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  5
        -----------
		Addr <=  "00000000000000";
		Trees_din <= x"05053e50";
		wait for Clk_period;
		Addr <=  "00000000000001";
		Trees_din <= x"05005828";
		wait for Clk_period;
		Addr <=  "00000000000010";
		Trees_din <= x"05fe4a0c";
		wait for Clk_period;
		Addr <=  "00000000000011";
		Trees_din <= x"0b074c04";
		wait for Clk_period;
		Addr <=  "00000000000100";
		Trees_din <= x"ff4e00b5";
		wait for Clk_period;
		Addr <=  "00000000000101";
		Trees_din <= x"05fd0e04";
		wait for Clk_period;
		Addr <=  "00000000000110";
		Trees_din <= x"ff6c00b5";
		wait for Clk_period;
		Addr <=  "00000000000111";
		Trees_din <= x"002700b5";
		wait for Clk_period;
		Addr <=  "00000000001000";
		Trees_din <= x"04001f0c";
		wait for Clk_period;
		Addr <=  "00000000001001";
		Trees_din <= x"00fce804";
		wait for Clk_period;
		Addr <=  "00000000001010";
		Trees_din <= x"005900b5";
		wait for Clk_period;
		Addr <=  "00000000001011";
		Trees_din <= x"0d000004";
		wait for Clk_period;
		Addr <=  "00000000001100";
		Trees_din <= x"fff100b5";
		wait for Clk_period;
		Addr <=  "00000000001101";
		Trees_din <= x"ff5100b5";
		wait for Clk_period;
		Addr <=  "00000000001110";
		Trees_din <= x"1403ab08";
		wait for Clk_period;
		Addr <=  "00000000001111";
		Trees_din <= x"19009204";
		wait for Clk_period;
		Addr <=  "00000000010000";
		Trees_din <= x"008900b5";
		wait for Clk_period;
		Addr <=  "00000000010001";
		Trees_din <= x"ff9a00b5";
		wait for Clk_period;
		Addr <=  "00000000010010";
		Trees_din <= x"13ffa004";
		wait for Clk_period;
		Addr <=  "00000000010011";
		Trees_din <= x"001200b5";
		wait for Clk_period;
		Addr <=  "00000000010100";
		Trees_din <= x"026000b5";
		wait for Clk_period;
		Addr <=  "00000000010101";
		Trees_din <= x"03fc2f18";
		wait for Clk_period;
		Addr <=  "00000000010110";
		Trees_din <= x"03fa9f0c";
		wait for Clk_period;
		Addr <=  "00000000010111";
		Trees_din <= x"1c002204";
		wait for Clk_period;
		Addr <=  "00000000011000";
		Trees_din <= x"ffe500b5";
		wait for Clk_period;
		Addr <=  "00000000011001";
		Trees_din <= x"0f000004";
		wait for Clk_period;
		Addr <=  "00000000011010";
		Trees_din <= x"ffda00b5";
		wait for Clk_period;
		Addr <=  "00000000011011";
		Trees_din <= x"ff5300b5";
		wait for Clk_period;
		Addr <=  "00000000011100";
		Trees_din <= x"05034408";
		wait for Clk_period;
		Addr <=  "00000000011101";
		Trees_din <= x"01ffb304";
		wait for Clk_period;
		Addr <=  "00000000011110";
		Trees_din <= x"ff6a00b5";
		wait for Clk_period;
		Addr <=  "00000000011111";
		Trees_din <= x"008e00b5";
		wait for Clk_period;
		Addr <=  "00000000100000";
		Trees_din <= x"013c00b5";
		wait for Clk_period;
		Addr <=  "00000000100001";
		Trees_din <= x"0208950c";
		wait for Clk_period;
		Addr <=  "00000000100010";
		Trees_din <= x"0009f008";
		wait for Clk_period;
		Addr <=  "00000000100011";
		Trees_din <= x"01011d04";
		wait for Clk_period;
		Addr <=  "00000000100100";
		Trees_din <= x"029700b5";
		wait for Clk_period;
		Addr <=  "00000000100101";
		Trees_din <= x"002700b5";
		wait for Clk_period;
		Addr <=  "00000000100110";
		Trees_din <= x"ff9d00b5";
		wait for Clk_period;
		Addr <=  "00000000100111";
		Trees_din <= x"ff8900b5";
		wait for Clk_period;
		Addr <=  "00000000101000";
		Trees_din <= x"06fb0208";
		wait for Clk_period;
		Addr <=  "00000000101001";
		Trees_din <= x"03f8a504";
		wait for Clk_period;
		Addr <=  "00000000101010";
		Trees_din <= x"ff7500b5";
		wait for Clk_period;
		Addr <=  "00000000101011";
		Trees_din <= x"00b200b5";
		wait for Clk_period;
		Addr <=  "00000000101100";
		Trees_din <= x"02b600b5";
		wait for Clk_period;
		Addr <=  "00000000101101";
		Trees_din <= x"05005840";
		wait for Clk_period;
		Addr <=  "00000000101110";
		Trees_din <= x"05fe4a14";
		wait for Clk_period;
		Addr <=  "00000000101111";
		Trees_din <= x"0b074c0c";
		wait for Clk_period;
		Addr <=  "00000000110000";
		Trees_din <= x"0a07cb04";
		wait for Clk_period;
		Addr <=  "00000000110001";
		Trees_din <= x"ff550199";
		wait for Clk_period;
		Addr <=  "00000000110010";
		Trees_din <= x"12003304";
		wait for Clk_period;
		Addr <=  "00000000110011";
		Trees_din <= x"ff740199";
		wait for Clk_period;
		Addr <=  "00000000110100";
		Trees_din <= x"00410199";
		wait for Clk_period;
		Addr <=  "00000000110101";
		Trees_din <= x"1b003b04";
		wait for Clk_period;
		Addr <=  "00000000110110";
		Trees_din <= x"ff760199";
		wait for Clk_period;
		Addr <=  "00000000110111";
		Trees_din <= x"003e0199";
		wait for Clk_period;
		Addr <=  "00000000111000";
		Trees_din <= x"04001f14";
		wait for Clk_period;
		Addr <=  "00000000111001";
		Trees_din <= x"00fce808";
		wait for Clk_period;
		Addr <=  "00000000111010";
		Trees_din <= x"0c00d004";
		wait for Clk_period;
		Addr <=  "00000000111011";
		Trees_din <= x"00d00199";
		wait for Clk_period;
		Addr <=  "00000000111100";
		Trees_din <= x"ffa40199";
		wait for Clk_period;
		Addr <=  "00000000111101";
		Trees_din <= x"0d000004";
		wait for Clk_period;
		Addr <=  "00000000111110";
		Trees_din <= x"ffff0199";
		wait for Clk_period;
		Addr <=  "00000000111111";
		Trees_din <= x"11fab304";
		wait for Clk_period;
		Addr <=  "00000001000000";
		Trees_din <= x"ffee0199";
		wait for Clk_period;
		Addr <=  "00000001000001";
		Trees_din <= x"ff570199";
		wait for Clk_period;
		Addr <=  "00000001000010";
		Trees_din <= x"1403ab10";
		wait for Clk_period;
		Addr <=  "00000001000011";
		Trees_din <= x"17020308";
		wait for Clk_period;
		Addr <=  "00000001000100";
		Trees_din <= x"14005904";
		wait for Clk_period;
		Addr <=  "00000001000101";
		Trees_din <= x"00ca0199";
		wait for Clk_period;
		Addr <=  "00000001000110";
		Trees_din <= x"ff800199";
		wait for Clk_period;
		Addr <=  "00000001000111";
		Trees_din <= x"1c002d04";
		wait for Clk_period;
		Addr <=  "00000001001000";
		Trees_din <= x"ffbb0199";
		wait for Clk_period;
		Addr <=  "00000001001001";
		Trees_din <= x"00ee0199";
		wait for Clk_period;
		Addr <=  "00000001001010";
		Trees_din <= x"1b003a04";
		wait for Clk_period;
		Addr <=  "00000001001011";
		Trees_din <= x"01850199";
		wait for Clk_period;
		Addr <=  "00000001001100";
		Trees_din <= x"000b0199";
		wait for Clk_period;
		Addr <=  "00000001001101";
		Trees_din <= x"000e4f24";
		wait for Clk_period;
		Addr <=  "00000001001110";
		Trees_din <= x"0209761c";
		wait for Clk_period;
		Addr <=  "00000001001111";
		Trees_din <= x"0501f810";
		wait for Clk_period;
		Addr <=  "00000001010000";
		Trees_din <= x"1004c508";
		wait for Clk_period;
		Addr <=  "00000001010001";
		Trees_din <= x"1600cd04";
		wait for Clk_period;
		Addr <=  "00000001010010";
		Trees_din <= x"ff800199";
		wait for Clk_period;
		Addr <=  "00000001010011";
		Trees_din <= x"01c80199";
		wait for Clk_period;
		Addr <=  "00000001010100";
		Trees_din <= x"06f84404";
		wait for Clk_period;
		Addr <=  "00000001010101";
		Trees_din <= x"00280199";
		wait for Clk_period;
		Addr <=  "00000001010110";
		Trees_din <= x"ff740199";
		wait for Clk_period;
		Addr <=  "00000001010111";
		Trees_din <= x"0b04c108";
		wait for Clk_period;
		Addr <=  "00000001011000";
		Trees_din <= x"07005c04";
		wait for Clk_period;
		Addr <=  "00000001011001";
		Trees_din <= x"02260199";
		wait for Clk_period;
		Addr <=  "00000001011010";
		Trees_din <= x"00ac0199";
		wait for Clk_period;
		Addr <=  "00000001011011";
		Trees_din <= x"008d0199";
		wait for Clk_period;
		Addr <=  "00000001011100";
		Trees_din <= x"06fbb604";
		wait for Clk_period;
		Addr <=  "00000001011101";
		Trees_din <= x"ff5e0199";
		wait for Clk_period;
		Addr <=  "00000001011110";
		Trees_din <= x"013b0199";
		wait for Clk_period;
		Addr <=  "00000001011111";
		Trees_din <= x"1c002204";
		wait for Clk_period;
		Addr <=  "00000001100000";
		Trees_din <= x"00020199";
		wait for Clk_period;
		Addr <=  "00000001100001";
		Trees_din <= x"0f000008";
		wait for Clk_period;
		Addr <=  "00000001100010";
		Trees_din <= x"03f4d804";
		wait for Clk_period;
		Addr <=  "00000001100011";
		Trees_din <= x"ffa50199";
		wait for Clk_period;
		Addr <=  "00000001100100";
		Trees_din <= x"00380199";
		wait for Clk_period;
		Addr <=  "00000001100101";
		Trees_din <= x"ff570199";
		wait for Clk_period;
		Addr <=  "00000001100110";
		Trees_din <= x"05005848";
		wait for Clk_period;
		Addr <=  "00000001100111";
		Trees_din <= x"05fe4a1c";
		wait for Clk_period;
		Addr <=  "00000001101000";
		Trees_din <= x"0b074c14";
		wait for Clk_period;
		Addr <=  "00000001101001";
		Trees_din <= x"0a07cb0c";
		wait for Clk_period;
		Addr <=  "00000001101010";
		Trees_din <= x"0e043204";
		wait for Clk_period;
		Addr <=  "00000001101011";
		Trees_din <= x"ff590275";
		wait for Clk_period;
		Addr <=  "00000001101100";
		Trees_din <= x"07004a04";
		wait for Clk_period;
		Addr <=  "00000001101101";
		Trees_din <= x"00a30275";
		wait for Clk_period;
		Addr <=  "00000001101110";
		Trees_din <= x"ff650275";
		wait for Clk_period;
		Addr <=  "00000001101111";
		Trees_din <= x"0e010504";
		wait for Clk_period;
		Addr <=  "00000001110000";
		Trees_din <= x"ff7c0275";
		wait for Clk_period;
		Addr <=  "00000001110001";
		Trees_din <= x"00420275";
		wait for Clk_period;
		Addr <=  "00000001110010";
		Trees_din <= x"15008d04";
		wait for Clk_period;
		Addr <=  "00000001110011";
		Trees_din <= x"00420275";
		wait for Clk_period;
		Addr <=  "00000001110100";
		Trees_din <= x"ff7e0275";
		wait for Clk_period;
		Addr <=  "00000001110101";
		Trees_din <= x"04001f14";
		wait for Clk_period;
		Addr <=  "00000001110110";
		Trees_din <= x"00fce808";
		wait for Clk_period;
		Addr <=  "00000001110111";
		Trees_din <= x"10041004";
		wait for Clk_period;
		Addr <=  "00000001111000";
		Trees_din <= x"ffa30275";
		wait for Clk_period;
		Addr <=  "00000001111001";
		Trees_din <= x"00c90275";
		wait for Clk_period;
		Addr <=  "00000001111010";
		Trees_din <= x"0d000004";
		wait for Clk_period;
		Addr <=  "00000001111011";
		Trees_din <= x"00080275";
		wait for Clk_period;
		Addr <=  "00000001111100";
		Trees_din <= x"11fab304";
		wait for Clk_period;
		Addr <=  "00000001111101";
		Trees_din <= x"fffa0275";
		wait for Clk_period;
		Addr <=  "00000001111110";
		Trees_din <= x"ff5c0275";
		wait for Clk_period;
		Addr <=  "00000001111111";
		Trees_din <= x"06f66f08";
		wait for Clk_period;
		Addr <=  "00000010000000";
		Trees_din <= x"09005b04";
		wait for Clk_period;
		Addr <=  "00000010000001";
		Trees_din <= x"ff620275";
		wait for Clk_period;
		Addr <=  "00000010000010";
		Trees_din <= x"00c80275";
		wait for Clk_period;
		Addr <=  "00000010000011";
		Trees_din <= x"01010a08";
		wait for Clk_period;
		Addr <=  "00000010000100";
		Trees_din <= x"09005304";
		wait for Clk_period;
		Addr <=  "00000010000101";
		Trees_din <= x"00930275";
		wait for Clk_period;
		Addr <=  "00000010000110";
		Trees_din <= x"ffa00275";
		wait for Clk_period;
		Addr <=  "00000010000111";
		Trees_din <= x"11025504";
		wait for Clk_period;
		Addr <=  "00000010001000";
		Trees_din <= x"01a40275";
		wait for Clk_period;
		Addr <=  "00000010001001";
		Trees_din <= x"00160275";
		wait for Clk_period;
		Addr <=  "00000010001010";
		Trees_din <= x"000e4f1c";
		wait for Clk_period;
		Addr <=  "00000010001011";
		Trees_din <= x"020c0718";
		wait for Clk_period;
		Addr <=  "00000010001100";
		Trees_din <= x"0501a40c";
		wait for Clk_period;
		Addr <=  "00000010001101";
		Trees_din <= x"10045108";
		wait for Clk_period;
		Addr <=  "00000010001110";
		Trees_din <= x"1600cd04";
		wait for Clk_period;
		Addr <=  "00000010001111";
		Trees_din <= x"ff800275";
		wait for Clk_period;
		Addr <=  "00000010010000";
		Trees_din <= x"01290275";
		wait for Clk_period;
		Addr <=  "00000010010001";
		Trees_din <= x"ff6f0275";
		wait for Clk_period;
		Addr <=  "00000010010010";
		Trees_din <= x"1f000008";
		wait for Clk_period;
		Addr <=  "00000010010011";
		Trees_din <= x"10f8a604";
		wait for Clk_period;
		Addr <=  "00000010010100";
		Trees_din <= x"00160275";
		wait for Clk_period;
		Addr <=  "00000010010101";
		Trees_din <= x"016b0275";
		wait for Clk_period;
		Addr <=  "00000010010110";
		Trees_din <= x"000b0275";
		wait for Clk_period;
		Addr <=  "00000010010111";
		Trees_din <= x"ff670275";
		wait for Clk_period;
		Addr <=  "00000010011000";
		Trees_din <= x"1c002204";
		wait for Clk_period;
		Addr <=  "00000010011001";
		Trees_din <= x"000c0275";
		wait for Clk_period;
		Addr <=  "00000010011010";
		Trees_din <= x"0f000004";
		wait for Clk_period;
		Addr <=  "00000010011011";
		Trees_din <= x"fff30275";
		wait for Clk_period;
		Addr <=  "00000010011100";
		Trees_din <= x"ff5c0275";
		wait for Clk_period;
		Addr <=  "00000010011101";
		Trees_din <= x"05005848";
		wait for Clk_period;
		Addr <=  "00000010011110";
		Trees_din <= x"05fe4a1c";
		wait for Clk_period;
		Addr <=  "00000010011111";
		Trees_din <= x"05fd3404";
		wait for Clk_period;
		Addr <=  "00000010100000";
		Trees_din <= x"ff5c0351";
		wait for Clk_period;
		Addr <=  "00000010100001";
		Trees_din <= x"0003e510";
		wait for Clk_period;
		Addr <=  "00000010100010";
		Trees_din <= x"09004a08";
		wait for Clk_period;
		Addr <=  "00000010100011";
		Trees_din <= x"0101c604";
		wait for Clk_period;
		Addr <=  "00000010100100";
		Trees_din <= x"001d0351";
		wait for Clk_period;
		Addr <=  "00000010100101";
		Trees_din <= x"016b0351";
		wait for Clk_period;
		Addr <=  "00000010100110";
		Trees_din <= x"11fd5b04";
		wait for Clk_period;
		Addr <=  "00000010100111";
		Trees_din <= x"00510351";
		wait for Clk_period;
		Addr <=  "00000010101000";
		Trees_din <= x"ff730351";
		wait for Clk_period;
		Addr <=  "00000010101001";
		Trees_din <= x"12047b04";
		wait for Clk_period;
		Addr <=  "00000010101010";
		Trees_din <= x"ff5d0351";
		wait for Clk_period;
		Addr <=  "00000010101011";
		Trees_din <= x"00290351";
		wait for Clk_period;
		Addr <=  "00000010101100";
		Trees_din <= x"03fbdc0c";
		wait for Clk_period;
		Addr <=  "00000010101101";
		Trees_din <= x"0d03d404";
		wait for Clk_period;
		Addr <=  "00000010101110";
		Trees_din <= x"ff5d0351";
		wait for Clk_period;
		Addr <=  "00000010101111";
		Trees_din <= x"15009504";
		wait for Clk_period;
		Addr <=  "00000010110000";
		Trees_din <= x"ff910351";
		wait for Clk_period;
		Addr <=  "00000010110001";
		Trees_din <= x"003e0351";
		wait for Clk_period;
		Addr <=  "00000010110010";
		Trees_din <= x"0c012a10";
		wait for Clk_period;
		Addr <=  "00000010110011";
		Trees_din <= x"08006608";
		wait for Clk_period;
		Addr <=  "00000010110100";
		Trees_din <= x"04070604";
		wait for Clk_period;
		Addr <=  "00000010110101";
		Trees_din <= x"ff6d0351";
		wait for Clk_period;
		Addr <=  "00000010110110";
		Trees_din <= x"00b50351";
		wait for Clk_period;
		Addr <=  "00000010110111";
		Trees_din <= x"18004904";
		wait for Clk_period;
		Addr <=  "00000010111000";
		Trees_din <= x"012a0351";
		wait for Clk_period;
		Addr <=  "00000010111001";
		Trees_din <= x"ff9a0351";
		wait for Clk_period;
		Addr <=  "00000010111010";
		Trees_din <= x"17000008";
		wait for Clk_period;
		Addr <=  "00000010111011";
		Trees_din <= x"11027004";
		wait for Clk_period;
		Addr <=  "00000010111100";
		Trees_din <= x"010a0351";
		wait for Clk_period;
		Addr <=  "00000010111101";
		Trees_din <= x"ff900351";
		wait for Clk_period;
		Addr <=  "00000010111110";
		Trees_din <= x"1400db04";
		wait for Clk_period;
		Addr <=  "00000010111111";
		Trees_din <= x"ffe80351";
		wait for Clk_period;
		Addr <=  "00000011000000";
		Trees_din <= x"ff5e0351";
		wait for Clk_period;
		Addr <=  "00000011000001";
		Trees_din <= x"000e4f1c";
		wait for Clk_period;
		Addr <=  "00000011000010";
		Trees_din <= x"020c0718";
		wait for Clk_period;
		Addr <=  "00000011000011";
		Trees_din <= x"0d03b210";
		wait for Clk_period;
		Addr <=  "00000011000100";
		Trees_din <= x"0501a408";
		wait for Clk_period;
		Addr <=  "00000011000101";
		Trees_din <= x"04fbe704";
		wait for Clk_period;
		Addr <=  "00000011000110";
		Trees_din <= x"ff750351";
		wait for Clk_period;
		Addr <=  "00000011000111";
		Trees_din <= x"00a60351";
		wait for Clk_period;
		Addr <=  "00000011001000";
		Trees_din <= x"0e045b04";
		wait for Clk_period;
		Addr <=  "00000011001001";
		Trees_din <= x"01270351";
		wait for Clk_period;
		Addr <=  "00000011001010";
		Trees_din <= x"fff50351";
		wait for Clk_period;
		Addr <=  "00000011001011";
		Trees_din <= x"08002d04";
		wait for Clk_period;
		Addr <=  "00000011001100";
		Trees_din <= x"ff950351";
		wait for Clk_period;
		Addr <=  "00000011001101";
		Trees_din <= x"00170351";
		wait for Clk_period;
		Addr <=  "00000011001110";
		Trees_din <= x"ff6d0351";
		wait for Clk_period;
		Addr <=  "00000011001111";
		Trees_din <= x"1c002204";
		wait for Clk_period;
		Addr <=  "00000011010000";
		Trees_din <= x"00160351";
		wait for Clk_period;
		Addr <=  "00000011010001";
		Trees_din <= x"020b0104";
		wait for Clk_period;
		Addr <=  "00000011010010";
		Trees_din <= x"ff600351";
		wait for Clk_period;
		Addr <=  "00000011010011";
		Trees_din <= x"00010351";
		wait for Clk_period;
		Addr <=  "00000011010100";
		Trees_din <= x"05005848";
		wait for Clk_period;
		Addr <=  "00000011010101";
		Trees_din <= x"05fe4a1c";
		wait for Clk_period;
		Addr <=  "00000011010110";
		Trees_din <= x"05fd3404";
		wait for Clk_period;
		Addr <=  "00000011010111";
		Trees_din <= x"ff5e041d";
		wait for Clk_period;
		Addr <=  "00000011011000";
		Trees_din <= x"0003e510";
		wait for Clk_period;
		Addr <=  "00000011011001";
		Trees_din <= x"09004a08";
		wait for Clk_period;
		Addr <=  "00000011011010";
		Trees_din <= x"09004504";
		wait for Clk_period;
		Addr <=  "00000011011011";
		Trees_din <= x"0006041d";
		wait for Clk_period;
		Addr <=  "00000011011100";
		Trees_din <= x"0167041d";
		wait for Clk_period;
		Addr <=  "00000011011101";
		Trees_din <= x"11fd5b04";
		wait for Clk_period;
		Addr <=  "00000011011110";
		Trees_din <= x"0049041d";
		wait for Clk_period;
		Addr <=  "00000011011111";
		Trees_din <= x"ff7a041d";
		wait for Clk_period;
		Addr <=  "00000011100000";
		Trees_din <= x"12047b04";
		wait for Clk_period;
		Addr <=  "00000011100001";
		Trees_din <= x"ff60041d";
		wait for Clk_period;
		Addr <=  "00000011100010";
		Trees_din <= x"002f041d";
		wait for Clk_period;
		Addr <=  "00000011100011";
		Trees_din <= x"03fbdc0c";
		wait for Clk_period;
		Addr <=  "00000011100100";
		Trees_din <= x"0d03d404";
		wait for Clk_period;
		Addr <=  "00000011100101";
		Trees_din <= x"ff60041d";
		wait for Clk_period;
		Addr <=  "00000011100110";
		Trees_din <= x"13ffa404";
		wait for Clk_period;
		Addr <=  "00000011100111";
		Trees_din <= x"ff99041d";
		wait for Clk_period;
		Addr <=  "00000011101000";
		Trees_din <= x"0044041d";
		wait for Clk_period;
		Addr <=  "00000011101001";
		Trees_din <= x"0c012a10";
		wait for Clk_period;
		Addr <=  "00000011101010";
		Trees_din <= x"08006608";
		wait for Clk_period;
		Addr <=  "00000011101011";
		Trees_din <= x"08000004";
		wait for Clk_period;
		Addr <=  "00000011101100";
		Trees_din <= x"00cb041d";
		wait for Clk_period;
		Addr <=  "00000011101101";
		Trees_din <= x"ff72041d";
		wait for Clk_period;
		Addr <=  "00000011101110";
		Trees_din <= x"09004d04";
		wait for Clk_period;
		Addr <=  "00000011101111";
		Trees_din <= x"ffcc041d";
		wait for Clk_period;
		Addr <=  "00000011110000";
		Trees_din <= x"0103041d";
		wait for Clk_period;
		Addr <=  "00000011110001";
		Trees_din <= x"17000008";
		wait for Clk_period;
		Addr <=  "00000011110010";
		Trees_din <= x"11027004";
		wait for Clk_period;
		Addr <=  "00000011110011";
		Trees_din <= x"00d1041d";
		wait for Clk_period;
		Addr <=  "00000011110100";
		Trees_din <= x"ff95041d";
		wait for Clk_period;
		Addr <=  "00000011110101";
		Trees_din <= x"1400db04";
		wait for Clk_period;
		Addr <=  "00000011110110";
		Trees_din <= x"fff0041d";
		wait for Clk_period;
		Addr <=  "00000011110111";
		Trees_din <= x"ff62041d";
		wait for Clk_period;
		Addr <=  "00000011111000";
		Trees_din <= x"000fd318";
		wait for Clk_period;
		Addr <=  "00000011111001";
		Trees_din <= x"020c0714";
		wait for Clk_period;
		Addr <=  "00000011111010";
		Trees_din <= x"06f53104";
		wait for Clk_period;
		Addr <=  "00000011111011";
		Trees_din <= x"ff89041d";
		wait for Clk_period;
		Addr <=  "00000011111100";
		Trees_din <= x"0d03b208";
		wait for Clk_period;
		Addr <=  "00000011111101";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00000011111110";
		Trees_din <= x"00de041d";
		wait for Clk_period;
		Addr <=  "00000011111111";
		Trees_din <= x"0047041d";
		wait for Clk_period;
		Addr <=  "00000100000000";
		Trees_din <= x"1b004504";
		wait for Clk_period;
		Addr <=  "00000100000001";
		Trees_din <= x"ff90041d";
		wait for Clk_period;
		Addr <=  "00000100000010";
		Trees_din <= x"0015041d";
		wait for Clk_period;
		Addr <=  "00000100000011";
		Trees_din <= x"ff73041d";
		wait for Clk_period;
		Addr <=  "00000100000100";
		Trees_din <= x"04fc4304";
		wait for Clk_period;
		Addr <=  "00000100000101";
		Trees_din <= x"ff63041d";
		wait for Clk_period;
		Addr <=  "00000100000110";
		Trees_din <= x"003f041d";
		wait for Clk_period;
		Addr <=  "00000100000111";
		Trees_din <= x"05005830";
		wait for Clk_period;
		Addr <=  "00000100001000";
		Trees_din <= x"05fd3404";
		wait for Clk_period;
		Addr <=  "00000100001001";
		Trees_din <= x"ff6004b9";
		wait for Clk_period;
		Addr <=  "00000100001010";
		Trees_din <= x"03fbdc10";
		wait for Clk_period;
		Addr <=  "00000100001011";
		Trees_din <= x"04fe1204";
		wait for Clk_period;
		Addr <=  "00000100001100";
		Trees_din <= x"ff6204b9";
		wait for Clk_period;
		Addr <=  "00000100001101";
		Trees_din <= x"0bfa8108";
		wait for Clk_period;
		Addr <=  "00000100001110";
		Trees_din <= x"06f5dc04";
		wait for Clk_period;
		Addr <=  "00000100001111";
		Trees_din <= x"00dc04b9";
		wait for Clk_period;
		Addr <=  "00000100010000";
		Trees_din <= x"ffac04b9";
		wait for Clk_period;
		Addr <=  "00000100010001";
		Trees_din <= x"ff7904b9";
		wait for Clk_period;
		Addr <=  "00000100010010";
		Trees_din <= x"0c012a10";
		wait for Clk_period;
		Addr <=  "00000100010011";
		Trees_din <= x"08006608";
		wait for Clk_period;
		Addr <=  "00000100010100";
		Trees_din <= x"08000004";
		wait for Clk_period;
		Addr <=  "00000100010101";
		Trees_din <= x"007704b9";
		wait for Clk_period;
		Addr <=  "00000100010110";
		Trees_din <= x"ff8e04b9";
		wait for Clk_period;
		Addr <=  "00000100010111";
		Trees_din <= x"0202b804";
		wait for Clk_period;
		Addr <=  "00000100011000";
		Trees_din <= x"00ad04b9";
		wait for Clk_period;
		Addr <=  "00000100011001";
		Trees_din <= x"ffca04b9";
		wait for Clk_period;
		Addr <=  "00000100011010";
		Trees_din <= x"0a04d608";
		wait for Clk_period;
		Addr <=  "00000100011011";
		Trees_din <= x"02fe7804";
		wait for Clk_period;
		Addr <=  "00000100011100";
		Trees_din <= x"fffb04b9";
		wait for Clk_period;
		Addr <=  "00000100011101";
		Trees_din <= x"ff7404b9";
		wait for Clk_period;
		Addr <=  "00000100011110";
		Trees_din <= x"009404b9";
		wait for Clk_period;
		Addr <=  "00000100011111";
		Trees_din <= x"03f79304";
		wait for Clk_period;
		Addr <=  "00000100100000";
		Trees_din <= x"ff6604b9";
		wait for Clk_period;
		Addr <=  "00000100100001";
		Trees_din <= x"020c0718";
		wait for Clk_period;
		Addr <=  "00000100100010";
		Trees_din <= x"000e4f10";
		wait for Clk_period;
		Addr <=  "00000100100011";
		Trees_din <= x"0501a408";
		wait for Clk_period;
		Addr <=  "00000100100100";
		Trees_din <= x"0801b804";
		wait for Clk_period;
		Addr <=  "00000100100101";
		Trees_din <= x"ffc504b9";
		wait for Clk_period;
		Addr <=  "00000100100110";
		Trees_din <= x"00a304b9";
		wait for Clk_period;
		Addr <=  "00000100100111";
		Trees_din <= x"0e045b04";
		wait for Clk_period;
		Addr <=  "00000100101000";
		Trees_din <= x"00d004b9";
		wait for Clk_period;
		Addr <=  "00000100101001";
		Trees_din <= x"ffe604b9";
		wait for Clk_period;
		Addr <=  "00000100101010";
		Trees_din <= x"08008f04";
		wait for Clk_period;
		Addr <=  "00000100101011";
		Trees_din <= x"008004b9";
		wait for Clk_period;
		Addr <=  "00000100101100";
		Trees_din <= x"ff7c04b9";
		wait for Clk_period;
		Addr <=  "00000100101101";
		Trees_din <= x"ff8104b9";
		wait for Clk_period;
		Addr <=  "00000100101110";
		Trees_din <= x"05fede2c";
		wait for Clk_period;
		Addr <=  "00000100101111";
		Trees_din <= x"05fd3404";
		wait for Clk_period;
		Addr <=  "00000100110000";
		Trees_din <= x"ff620575";
		wait for Clk_period;
		Addr <=  "00000100110001";
		Trees_din <= x"04065f18";
		wait for Clk_period;
		Addr <=  "00000100110010";
		Trees_din <= x"0e043210";
		wait for Clk_period;
		Addr <=  "00000100110011";
		Trees_din <= x"0104a608";
		wait for Clk_period;
		Addr <=  "00000100110100";
		Trees_din <= x"16000604";
		wait for Clk_period;
		Addr <=  "00000100110101";
		Trees_din <= x"ffce0575";
		wait for Clk_period;
		Addr <=  "00000100110110";
		Trees_din <= x"ff610575";
		wait for Clk_period;
		Addr <=  "00000100110111";
		Trees_din <= x"1603f904";
		wait for Clk_period;
		Addr <=  "00000100111000";
		Trees_din <= x"ff830575";
		wait for Clk_period;
		Addr <=  "00000100111001";
		Trees_din <= x"008f0575";
		wait for Clk_period;
		Addr <=  "00000100111010";
		Trees_din <= x"000d9f04";
		wait for Clk_period;
		Addr <=  "00000100111011";
		Trees_din <= x"00e30575";
		wait for Clk_period;
		Addr <=  "00000100111100";
		Trees_din <= x"ff880575";
		wait for Clk_period;
		Addr <=  "00000100111101";
		Trees_din <= x"18004308";
		wait for Clk_period;
		Addr <=  "00000100111110";
		Trees_din <= x"1c002804";
		wait for Clk_period;
		Addr <=  "00000100111111";
		Trees_din <= x"00150575";
		wait for Clk_period;
		Addr <=  "00000101000000";
		Trees_din <= x"ff7e0575";
		wait for Clk_period;
		Addr <=  "00000101000001";
		Trees_din <= x"06f76004";
		wait for Clk_period;
		Addr <=  "00000101000010";
		Trees_din <= x"01410575";
		wait for Clk_period;
		Addr <=  "00000101000011";
		Trees_din <= x"ff940575";
		wait for Clk_period;
		Addr <=  "00000101000100";
		Trees_din <= x"0009f01c";
		wait for Clk_period;
		Addr <=  "00000101000101";
		Trees_din <= x"02097614";
		wait for Clk_period;
		Addr <=  "00000101000110";
		Trees_din <= x"0d03530c";
		wait for Clk_period;
		Addr <=  "00000101000111";
		Trees_din <= x"06f55c04";
		wait for Clk_period;
		Addr <=  "00000101001000";
		Trees_din <= x"ff8f0575";
		wait for Clk_period;
		Addr <=  "00000101001001";
		Trees_din <= x"12028704";
		wait for Clk_period;
		Addr <=  "00000101001010";
		Trees_din <= x"00a50575";
		wait for Clk_period;
		Addr <=  "00000101001011";
		Trees_din <= x"00030575";
		wait for Clk_period;
		Addr <=  "00000101001100";
		Trees_din <= x"02fe6f04";
		wait for Clk_period;
		Addr <=  "00000101001101";
		Trees_din <= x"00630575";
		wait for Clk_period;
		Addr <=  "00000101001110";
		Trees_din <= x"ff790575";
		wait for Clk_period;
		Addr <=  "00000101001111";
		Trees_din <= x"06fbb604";
		wait for Clk_period;
		Addr <=  "00000101010000";
		Trees_din <= x"ff6d0575";
		wait for Clk_period;
		Addr <=  "00000101010001";
		Trees_din <= x"009d0575";
		wait for Clk_period;
		Addr <=  "00000101010010";
		Trees_din <= x"06f9ff0c";
		wait for Clk_period;
		Addr <=  "00000101010011";
		Trees_din <= x"0b069b08";
		wait for Clk_period;
		Addr <=  "00000101010100";
		Trees_din <= x"0f000004";
		wait for Clk_period;
		Addr <=  "00000101010101";
		Trees_din <= x"00130575";
		wait for Clk_period;
		Addr <=  "00000101010110";
		Trees_din <= x"ff630575";
		wait for Clk_period;
		Addr <=  "00000101010111";
		Trees_din <= x"001c0575";
		wait for Clk_period;
		Addr <=  "00000101011000";
		Trees_din <= x"000e4f04";
		wait for Clk_period;
		Addr <=  "00000101011001";
		Trees_din <= x"00ad0575";
		wait for Clk_period;
		Addr <=  "00000101011010";
		Trees_din <= x"09004c04";
		wait for Clk_period;
		Addr <=  "00000101011011";
		Trees_din <= x"00420575";
		wait for Clk_period;
		Addr <=  "00000101011100";
		Trees_din <= x"ff7a0575";
		wait for Clk_period;
		Addr <=  "00000101011101";
		Trees_din <= x"05fede30";
		wait for Clk_period;
		Addr <=  "00000101011110";
		Trees_din <= x"05fd3404";
		wait for Clk_period;
		Addr <=  "00000101011111";
		Trees_din <= x"ff630629";
		wait for Clk_period;
		Addr <=  "00000101100000";
		Trees_din <= x"04065f18";
		wait for Clk_period;
		Addr <=  "00000101100001";
		Trees_din <= x"0e043210";
		wait for Clk_period;
		Addr <=  "00000101100010";
		Trees_din <= x"0bfa2308";
		wait for Clk_period;
		Addr <=  "00000101100011";
		Trees_din <= x"04fe1204";
		wait for Clk_period;
		Addr <=  "00000101100100";
		Trees_din <= x"ff700629";
		wait for Clk_period;
		Addr <=  "00000101100101";
		Trees_din <= x"00430629";
		wait for Clk_period;
		Addr <=  "00000101100110";
		Trees_din <= x"1500b304";
		wait for Clk_period;
		Addr <=  "00000101100111";
		Trees_din <= x"ff620629";
		wait for Clk_period;
		Addr <=  "00000101101000";
		Trees_din <= x"001a0629";
		wait for Clk_period;
		Addr <=  "00000101101001";
		Trees_din <= x"000d9f04";
		wait for Clk_period;
		Addr <=  "00000101101010";
		Trees_din <= x"00c20629";
		wait for Clk_period;
		Addr <=  "00000101101011";
		Trees_din <= x"ff8f0629";
		wait for Clk_period;
		Addr <=  "00000101101100";
		Trees_din <= x"02fd8d04";
		wait for Clk_period;
		Addr <=  "00000101101101";
		Trees_din <= x"ff810629";
		wait for Clk_period;
		Addr <=  "00000101101110";
		Trees_din <= x"18004308";
		wait for Clk_period;
		Addr <=  "00000101101111";
		Trees_din <= x"0f03ba04";
		wait for Clk_period;
		Addr <=  "00000101110000";
		Trees_din <= x"ff9e0629";
		wait for Clk_period;
		Addr <=  "00000101110001";
		Trees_din <= x"00160629";
		wait for Clk_period;
		Addr <=  "00000101110010";
		Trees_din <= x"00fe2904";
		wait for Clk_period;
		Addr <=  "00000101110011";
		Trees_din <= x"013b0629";
		wait for Clk_period;
		Addr <=  "00000101110100";
		Trees_din <= x"00190629";
		wait for Clk_period;
		Addr <=  "00000101110101";
		Trees_din <= x"000fd324";
		wait for Clk_period;
		Addr <=  "00000101110110";
		Trees_din <= x"020c0720";
		wait for Clk_period;
		Addr <=  "00000101110111";
		Trees_din <= x"05024c10";
		wait for Clk_period;
		Addr <=  "00000101111000";
		Trees_din <= x"11fea808";
		wait for Clk_period;
		Addr <=  "00000101111001";
		Trees_din <= x"01005e04";
		wait for Clk_period;
		Addr <=  "00000101111010";
		Trees_din <= x"00ec0629";
		wait for Clk_period;
		Addr <=  "00000101111011";
		Trees_din <= x"fffd0629";
		wait for Clk_period;
		Addr <=  "00000101111100";
		Trees_din <= x"04fd5304";
		wait for Clk_period;
		Addr <=  "00000101111101";
		Trees_din <= x"ff860629";
		wait for Clk_period;
		Addr <=  "00000101111110";
		Trees_din <= x"00250629";
		wait for Clk_period;
		Addr <=  "00000101111111";
		Trees_din <= x"06f76008";
		wait for Clk_period;
		Addr <=  "00000110000000";
		Trees_din <= x"0afad104";
		wait for Clk_period;
		Addr <=  "00000110000001";
		Trees_din <= x"005d0629";
		wait for Clk_period;
		Addr <=  "00000110000010";
		Trees_din <= x"ff9f0629";
		wait for Clk_period;
		Addr <=  "00000110000011";
		Trees_din <= x"07005c04";
		wait for Clk_period;
		Addr <=  "00000110000100";
		Trees_din <= x"00b80629";
		wait for Clk_period;
		Addr <=  "00000110000101";
		Trees_din <= x"fff50629";
		wait for Clk_period;
		Addr <=  "00000110000110";
		Trees_din <= x"ff770629";
		wait for Clk_period;
		Addr <=  "00000110000111";
		Trees_din <= x"1c002204";
		wait for Clk_period;
		Addr <=  "00000110001000";
		Trees_din <= x"00210629";
		wait for Clk_period;
		Addr <=  "00000110001001";
		Trees_din <= x"ff680629";
		wait for Clk_period;
		Addr <=  "00000110001010";
		Trees_din <= x"05fe4a28";
		wait for Clk_period;
		Addr <=  "00000110001011";
		Trees_din <= x"05fd340c";
		wait for Clk_period;
		Addr <=  "00000110001100";
		Trees_din <= x"02fc0c08";
		wait for Clk_period;
		Addr <=  "00000110001101";
		Trees_din <= x"0e03b204";
		wait for Clk_period;
		Addr <=  "00000110001110";
		Trees_din <= x"ff7c06bd";
		wait for Clk_period;
		Addr <=  "00000110001111";
		Trees_din <= x"004506bd";
		wait for Clk_period;
		Addr <=  "00000110010000";
		Trees_din <= x"ff6306bd";
		wait for Clk_period;
		Addr <=  "00000110010001";
		Trees_din <= x"0003e514";
		wait for Clk_period;
		Addr <=  "00000110010010";
		Trees_din <= x"17004d04";
		wait for Clk_period;
		Addr <=  "00000110010011";
		Trees_din <= x"ff7506bd";
		wait for Clk_period;
		Addr <=  "00000110010100";
		Trees_din <= x"00025708";
		wait for Clk_period;
		Addr <=  "00000110010101";
		Trees_din <= x"04077804";
		wait for Clk_period;
		Addr <=  "00000110010110";
		Trees_din <= x"ff8306bd";
		wait for Clk_period;
		Addr <=  "00000110010111";
		Trees_din <= x"007706bd";
		wait for Clk_period;
		Addr <=  "00000110011000";
		Trees_din <= x"1004bf04";
		wait for Clk_period;
		Addr <=  "00000110011001";
		Trees_din <= x"015906bd";
		wait for Clk_period;
		Addr <=  "00000110011010";
		Trees_din <= x"003206bd";
		wait for Clk_period;
		Addr <=  "00000110011011";
		Trees_din <= x"1301d604";
		wait for Clk_period;
		Addr <=  "00000110011100";
		Trees_din <= x"ff6806bd";
		wait for Clk_period;
		Addr <=  "00000110011101";
		Trees_din <= x"002f06bd";
		wait for Clk_period;
		Addr <=  "00000110011110";
		Trees_din <= x"000fd31c";
		wait for Clk_period;
		Addr <=  "00000110011111";
		Trees_din <= x"06f56504";
		wait for Clk_period;
		Addr <=  "00000110100000";
		Trees_din <= x"ff6f06bd";
		wait for Clk_period;
		Addr <=  "00000110100001";
		Trees_din <= x"11043c10";
		wait for Clk_period;
		Addr <=  "00000110100010";
		Trees_din <= x"0e025f08";
		wait for Clk_period;
		Addr <=  "00000110100011";
		Trees_din <= x"0d038c04";
		wait for Clk_period;
		Addr <=  "00000110100100";
		Trees_din <= x"003506bd";
		wait for Clk_period;
		Addr <=  "00000110100101";
		Trees_din <= x"ff9006bd";
		wait for Clk_period;
		Addr <=  "00000110100110";
		Trees_din <= x"1203f704";
		wait for Clk_period;
		Addr <=  "00000110100111";
		Trees_din <= x"00c506bd";
		wait for Clk_period;
		Addr <=  "00000110101000";
		Trees_din <= x"000706bd";
		wait for Clk_period;
		Addr <=  "00000110101001";
		Trees_din <= x"09005704";
		wait for Clk_period;
		Addr <=  "00000110101010";
		Trees_din <= x"ff6406bd";
		wait for Clk_period;
		Addr <=  "00000110101011";
		Trees_din <= x"005c06bd";
		wait for Clk_period;
		Addr <=  "00000110101100";
		Trees_din <= x"1c002204";
		wait for Clk_period;
		Addr <=  "00000110101101";
		Trees_din <= x"000306bd";
		wait for Clk_period;
		Addr <=  "00000110101110";
		Trees_din <= x"ff6806bd";
		wait for Clk_period;
		Addr <=  "00000110101111";
		Trees_din <= x"05fe4a28";
		wait for Clk_period;
		Addr <=  "00000110110000";
		Trees_din <= x"05fd340c";
		wait for Clk_period;
		Addr <=  "00000110110001";
		Trees_din <= x"02fc0c08";
		wait for Clk_period;
		Addr <=  "00000110110010";
		Trees_din <= x"02fbdf04";
		wait for Clk_period;
		Addr <=  "00000110110011";
		Trees_din <= x"ff810759";
		wait for Clk_period;
		Addr <=  "00000110110100";
		Trees_din <= x"00490759";
		wait for Clk_period;
		Addr <=  "00000110110101";
		Trees_din <= x"ff640759";
		wait for Clk_period;
		Addr <=  "00000110110110";
		Trees_din <= x"0003e514";
		wait for Clk_period;
		Addr <=  "00000110110111";
		Trees_din <= x"17004d04";
		wait for Clk_period;
		Addr <=  "00000110111000";
		Trees_din <= x"ff790759";
		wait for Clk_period;
		Addr <=  "00000110111001";
		Trees_din <= x"00025708";
		wait for Clk_period;
		Addr <=  "00000110111010";
		Trees_din <= x"1300d304";
		wait for Clk_period;
		Addr <=  "00000110111011";
		Trees_din <= x"ffab0759";
		wait for Clk_period;
		Addr <=  "00000110111100";
		Trees_din <= x"00b10759";
		wait for Clk_period;
		Addr <=  "00000110111101";
		Trees_din <= x"03fe5104";
		wait for Clk_period;
		Addr <=  "00000110111110";
		Trees_din <= x"001e0759";
		wait for Clk_period;
		Addr <=  "00000110111111";
		Trees_din <= x"01410759";
		wait for Clk_period;
		Addr <=  "00000111000000";
		Trees_din <= x"1301d604";
		wait for Clk_period;
		Addr <=  "00000111000001";
		Trees_din <= x"ff6a0759";
		wait for Clk_period;
		Addr <=  "00000111000010";
		Trees_din <= x"00310759";
		wait for Clk_period;
		Addr <=  "00000111000011";
		Trees_din <= x"000fd320";
		wait for Clk_period;
		Addr <=  "00000111000100";
		Trees_din <= x"06f56504";
		wait for Clk_period;
		Addr <=  "00000111000101";
		Trees_din <= x"ff740759";
		wait for Clk_period;
		Addr <=  "00000111000110";
		Trees_din <= x"0502b810";
		wait for Clk_period;
		Addr <=  "00000111000111";
		Trees_din <= x"04fd2008";
		wait for Clk_period;
		Addr <=  "00000111001000";
		Trees_din <= x"1b004504";
		wait for Clk_period;
		Addr <=  "00000111001001";
		Trees_din <= x"ff6e0759";
		wait for Clk_period;
		Addr <=  "00000111001010";
		Trees_din <= x"008a0759";
		wait for Clk_period;
		Addr <=  "00000111001011";
		Trees_din <= x"0c010704";
		wait for Clk_period;
		Addr <=  "00000111001100";
		Trees_din <= x"007e0759";
		wait for Clk_period;
		Addr <=  "00000111001101";
		Trees_din <= x"00050759";
		wait for Clk_period;
		Addr <=  "00000111001110";
		Trees_din <= x"1103e208";
		wait for Clk_period;
		Addr <=  "00000111001111";
		Trees_din <= x"06f6f104";
		wait for Clk_period;
		Addr <=  "00000111010000";
		Trees_din <= x"fff30759";
		wait for Clk_period;
		Addr <=  "00000111010001";
		Trees_din <= x"00a30759";
		wait for Clk_period;
		Addr <=  "00000111010010";
		Trees_din <= x"ffcb0759";
		wait for Clk_period;
		Addr <=  "00000111010011";
		Trees_din <= x"1900b004";
		wait for Clk_period;
		Addr <=  "00000111010100";
		Trees_din <= x"ff6a0759";
		wait for Clk_period;
		Addr <=  "00000111010101";
		Trees_din <= x"00110759";
		wait for Clk_period;
		Addr <=  "00000111010110";
		Trees_din <= x"05fe4a28";
		wait for Clk_period;
		Addr <=  "00000111010111";
		Trees_din <= x"05fd340c";
		wait for Clk_period;
		Addr <=  "00000111011000";
		Trees_din <= x"02fc0c08";
		wait for Clk_period;
		Addr <=  "00000111011001";
		Trees_din <= x"02fbdf04";
		wait for Clk_period;
		Addr <=  "00000111011010";
		Trees_din <= x"ff8707f5";
		wait for Clk_period;
		Addr <=  "00000111011011";
		Trees_din <= x"004907f5";
		wait for Clk_period;
		Addr <=  "00000111011100";
		Trees_din <= x"ff6507f5";
		wait for Clk_period;
		Addr <=  "00000111011101";
		Trees_din <= x"0e043214";
		wait for Clk_period;
		Addr <=  "00000111011110";
		Trees_din <= x"1500b310";
		wait for Clk_period;
		Addr <=  "00000111011111";
		Trees_din <= x"1301c408";
		wait for Clk_period;
		Addr <=  "00000111100000";
		Trees_din <= x"02fd2b04";
		wait for Clk_period;
		Addr <=  "00000111100001";
		Trees_din <= x"ffe107f5";
		wait for Clk_period;
		Addr <=  "00000111100010";
		Trees_din <= x"ff6907f5";
		wait for Clk_period;
		Addr <=  "00000111100011";
		Trees_din <= x"00fe2904";
		wait for Clk_period;
		Addr <=  "00000111100100";
		Trees_din <= x"009f07f5";
		wait for Clk_period;
		Addr <=  "00000111100101";
		Trees_din <= x"ffa407f5";
		wait for Clk_period;
		Addr <=  "00000111100110";
		Trees_din <= x"004c07f5";
		wait for Clk_period;
		Addr <=  "00000111100111";
		Trees_din <= x"01060b04";
		wait for Clk_period;
		Addr <=  "00000111101000";
		Trees_din <= x"fff207f5";
		wait for Clk_period;
		Addr <=  "00000111101001";
		Trees_din <= x"00c507f5";
		wait for Clk_period;
		Addr <=  "00000111101010";
		Trees_din <= x"03f7a104";
		wait for Clk_period;
		Addr <=  "00000111101011";
		Trees_din <= x"ff6c07f5";
		wait for Clk_period;
		Addr <=  "00000111101100";
		Trees_din <= x"06f56504";
		wait for Clk_period;
		Addr <=  "00000111101101";
		Trees_din <= x"ff7b07f5";
		wait for Clk_period;
		Addr <=  "00000111101110";
		Trees_din <= x"12fea810";
		wait for Clk_period;
		Addr <=  "00000111101111";
		Trees_din <= x"07005708";
		wait for Clk_period;
		Addr <=  "00000111110000";
		Trees_din <= x"02ff3c04";
		wait for Clk_period;
		Addr <=  "00000111110001";
		Trees_din <= x"002207f5";
		wait for Clk_period;
		Addr <=  "00000111110010";
		Trees_din <= x"00d407f5";
		wait for Clk_period;
		Addr <=  "00000111110011";
		Trees_din <= x"1d004404";
		wait for Clk_period;
		Addr <=  "00000111110100";
		Trees_din <= x"ff8d07f5";
		wait for Clk_period;
		Addr <=  "00000111110101";
		Trees_din <= x"006107f5";
		wait for Clk_period;
		Addr <=  "00000111110110";
		Trees_din <= x"01038908";
		wait for Clk_period;
		Addr <=  "00000111110111";
		Trees_din <= x"0500f004";
		wait for Clk_period;
		Addr <=  "00000111111000";
		Trees_din <= x"ffd107f5";
		wait for Clk_period;
		Addr <=  "00000111111001";
		Trees_din <= x"004307f5";
		wait for Clk_period;
		Addr <=  "00000111111010";
		Trees_din <= x"0a024104";
		wait for Clk_period;
		Addr <=  "00000111111011";
		Trees_din <= x"000e07f5";
		wait for Clk_period;
		Addr <=  "00000111111100";
		Trees_din <= x"012a07f5";
		wait for Clk_period;
		Addr <=  "00000111111101";
		Trees_din <= x"05fd4e14";
		wait for Clk_period;
		Addr <=  "00000111111110";
		Trees_din <= x"02fc0c08";
		wait for Clk_period;
		Addr <=  "00000111111111";
		Trees_din <= x"0103e604";
		wait for Clk_period;
		Addr <=  "00001000000000";
		Trees_din <= x"ff8c0871";
		wait for Clk_period;
		Addr <=  "00001000000001";
		Trees_din <= x"00490871";
		wait for Clk_period;
		Addr <=  "00001000000010";
		Trees_din <= x"05fd3404";
		wait for Clk_period;
		Addr <=  "00001000000011";
		Trees_din <= x"ff660871";
		wait for Clk_period;
		Addr <=  "00001000000100";
		Trees_din <= x"0f02fb04";
		wait for Clk_period;
		Addr <=  "00001000000101";
		Trees_din <= x"ff920871";
		wait for Clk_period;
		Addr <=  "00001000000110";
		Trees_din <= x"00210871";
		wait for Clk_period;
		Addr <=  "00001000000111";
		Trees_din <= x"000fd324";
		wait for Clk_period;
		Addr <=  "00001000001000";
		Trees_din <= x"06f50204";
		wait for Clk_period;
		Addr <=  "00001000001001";
		Trees_din <= x"ff760871";
		wait for Clk_period;
		Addr <=  "00001000001010";
		Trees_din <= x"01038910";
		wait for Clk_period;
		Addr <=  "00001000001011";
		Trees_din <= x"05005808";
		wait for Clk_period;
		Addr <=  "00001000001100";
		Trees_din <= x"02031004";
		wait for Clk_period;
		Addr <=  "00001000001101";
		Trees_din <= x"000d0871";
		wait for Clk_period;
		Addr <=  "00001000001110";
		Trees_din <= x"ff6c0871";
		wait for Clk_period;
		Addr <=  "00001000001111";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00001000010000";
		Trees_din <= x"00600871";
		wait for Clk_period;
		Addr <=  "00001000010001";
		Trees_din <= x"fff20871";
		wait for Clk_period;
		Addr <=  "00001000010010";
		Trees_din <= x"0c008c08";
		wait for Clk_period;
		Addr <=  "00001000010011";
		Trees_din <= x"0c004104";
		wait for Clk_period;
		Addr <=  "00001000010100";
		Trees_din <= x"002a0871";
		wait for Clk_period;
		Addr <=  "00001000010101";
		Trees_din <= x"014e0871";
		wait for Clk_period;
		Addr <=  "00001000010110";
		Trees_din <= x"00058404";
		wait for Clk_period;
		Addr <=  "00001000010111";
		Trees_din <= x"00800871";
		wait for Clk_period;
		Addr <=  "00001000011000";
		Trees_din <= x"ff850871";
		wait for Clk_period;
		Addr <=  "00001000011001";
		Trees_din <= x"1900b004";
		wait for Clk_period;
		Addr <=  "00001000011010";
		Trees_din <= x"ff6b0871";
		wait for Clk_period;
		Addr <=  "00001000011011";
		Trees_din <= x"00120871";
		wait for Clk_period;
		Addr <=  "00001000011100";
		Trees_din <= x"05fd4e14";
		wait for Clk_period;
		Addr <=  "00001000011101";
		Trees_din <= x"1104aa0c";
		wait for Clk_period;
		Addr <=  "00001000011110";
		Trees_din <= x"05fd3404";
		wait for Clk_period;
		Addr <=  "00001000011111";
		Trees_din <= x"ff6608e5";
		wait for Clk_period;
		Addr <=  "00001000100000";
		Trees_din <= x"0f02fb04";
		wait for Clk_period;
		Addr <=  "00001000100001";
		Trees_din <= x"ff9b08e5";
		wait for Clk_period;
		Addr <=  "00001000100010";
		Trees_din <= x"001c08e5";
		wait for Clk_period;
		Addr <=  "00001000100011";
		Trees_din <= x"04014904";
		wait for Clk_period;
		Addr <=  "00001000100100";
		Trees_din <= x"ff9308e5";
		wait for Clk_period;
		Addr <=  "00001000100101";
		Trees_din <= x"004608e5";
		wait for Clk_period;
		Addr <=  "00001000100110";
		Trees_din <= x"03f7a104";
		wait for Clk_period;
		Addr <=  "00001000100111";
		Trees_din <= x"ff6e08e5";
		wait for Clk_period;
		Addr <=  "00001000101000";
		Trees_din <= x"06f50204";
		wait for Clk_period;
		Addr <=  "00001000101001";
		Trees_din <= x"ff7c08e5";
		wait for Clk_period;
		Addr <=  "00001000101010";
		Trees_din <= x"07005810";
		wait for Clk_period;
		Addr <=  "00001000101011";
		Trees_din <= x"07005508";
		wait for Clk_period;
		Addr <=  "00001000101100";
		Trees_din <= x"00090504";
		wait for Clk_period;
		Addr <=  "00001000101101";
		Trees_din <= x"001708e5";
		wait for Clk_period;
		Addr <=  "00001000101110";
		Trees_din <= x"ff7a08e5";
		wait for Clk_period;
		Addr <=  "00001000101111";
		Trees_din <= x"0c023104";
		wait for Clk_period;
		Addr <=  "00001000110000";
		Trees_din <= x"00a608e5";
		wait for Clk_period;
		Addr <=  "00001000110001";
		Trees_din <= x"ffea08e5";
		wait for Clk_period;
		Addr <=  "00001000110010";
		Trees_din <= x"1301ab08";
		wait for Clk_period;
		Addr <=  "00001000110011";
		Trees_din <= x"1702c804";
		wait for Clk_period;
		Addr <=  "00001000110100";
		Trees_din <= x"ffb608e5";
		wait for Clk_period;
		Addr <=  "00001000110101";
		Trees_din <= x"002c08e5";
		wait for Clk_period;
		Addr <=  "00001000110110";
		Trees_din <= x"0afd2a04";
		wait for Clk_period;
		Addr <=  "00001000110111";
		Trees_din <= x"00b508e5";
		wait for Clk_period;
		Addr <=  "00001000111000";
		Trees_din <= x"002108e5";
		wait for Clk_period;
		Addr <=  "00001000111001";
		Trees_din <= x"05fd340c";
		wait for Clk_period;
		Addr <=  "00001000111010";
		Trees_din <= x"02fc0c08";
		wait for Clk_period;
		Addr <=  "00001000111011";
		Trees_din <= x"17000104";
		wait for Clk_period;
		Addr <=  "00001000111100";
		Trees_din <= x"00450981";
		wait for Clk_period;
		Addr <=  "00001000111101";
		Trees_din <= x"ff9d0981";
		wait for Clk_period;
		Addr <=  "00001000111110";
		Trees_din <= x"ff670981";
		wait for Clk_period;
		Addr <=  "00001000111111";
		Trees_din <= x"03f7a104";
		wait for Clk_period;
		Addr <=  "00001001000000";
		Trees_din <= x"ff700981";
		wait for Clk_period;
		Addr <=  "00001001000001";
		Trees_din <= x"05005820";
		wait for Clk_period;
		Addr <=  "00001001000010";
		Trees_din <= x"13fe5a10";
		wait for Clk_period;
		Addr <=  "00001001000011";
		Trees_din <= x"1500ae08";
		wait for Clk_period;
		Addr <=  "00001001000100";
		Trees_din <= x"04065f04";
		wait for Clk_period;
		Addr <=  "00001001000101";
		Trees_din <= x"ff770981";
		wait for Clk_period;
		Addr <=  "00001001000110";
		Trees_din <= x"00280981";
		wait for Clk_period;
		Addr <=  "00001001000111";
		Trees_din <= x"0af7d004";
		wait for Clk_period;
		Addr <=  "00001001001000";
		Trees_din <= x"00b10981";
		wait for Clk_period;
		Addr <=  "00001001001001";
		Trees_din <= x"000e0981";
		wait for Clk_period;
		Addr <=  "00001001001010";
		Trees_din <= x"1b003c08";
		wait for Clk_period;
		Addr <=  "00001001001011";
		Trees_din <= x"1400fa04";
		wait for Clk_period;
		Addr <=  "00001001001100";
		Trees_din <= x"00a10981";
		wait for Clk_period;
		Addr <=  "00001001001101";
		Trees_din <= x"fffb0981";
		wait for Clk_period;
		Addr <=  "00001001001110";
		Trees_din <= x"0b064804";
		wait for Clk_period;
		Addr <=  "00001001001111";
		Trees_din <= x"ff6f0981";
		wait for Clk_period;
		Addr <=  "00001001010000";
		Trees_din <= x"00a30981";
		wait for Clk_period;
		Addr <=  "00001001010001";
		Trees_din <= x"20040010";
		wait for Clk_period;
		Addr <=  "00001001010010";
		Trees_din <= x"1a00d308";
		wait for Clk_period;
		Addr <=  "00001001010011";
		Trees_din <= x"0f02a004";
		wait for Clk_period;
		Addr <=  "00001001010100";
		Trees_din <= x"ff680981";
		wait for Clk_period;
		Addr <=  "00001001010101";
		Trees_din <= x"002e0981";
		wait for Clk_period;
		Addr <=  "00001001010110";
		Trees_din <= x"0c014c04";
		wait for Clk_period;
		Addr <=  "00001001010111";
		Trees_din <= x"007a0981";
		wait for Clk_period;
		Addr <=  "00001001011000";
		Trees_din <= x"ffe60981";
		wait for Clk_period;
		Addr <=  "00001001011001";
		Trees_din <= x"1600db08";
		wait for Clk_period;
		Addr <=  "00001001011010";
		Trees_din <= x"0501f804";
		wait for Clk_period;
		Addr <=  "00001001011011";
		Trees_din <= x"ff7e0981";
		wait for Clk_period;
		Addr <=  "00001001011100";
		Trees_din <= x"00680981";
		wait for Clk_period;
		Addr <=  "00001001011101";
		Trees_din <= x"0c00b304";
		wait for Clk_period;
		Addr <=  "00001001011110";
		Trees_din <= x"ffda0981";
		wait for Clk_period;
		Addr <=  "00001001011111";
		Trees_din <= x"00970981";
		wait for Clk_period;
		Addr <=  "00001001100000";
		Trees_din <= x"05fd340c";
		wait for Clk_period;
		Addr <=  "00001001100001";
		Trees_din <= x"1104aa04";
		wait for Clk_period;
		Addr <=  "00001001100010";
		Trees_din <= x"ff6709e5";
		wait for Clk_period;
		Addr <=  "00001001100011";
		Trees_din <= x"0c02ca04";
		wait for Clk_period;
		Addr <=  "00001001100100";
		Trees_din <= x"ffa409e5";
		wait for Clk_period;
		Addr <=  "00001001100101";
		Trees_din <= x"004509e5";
		wait for Clk_period;
		Addr <=  "00001001100110";
		Trees_din <= x"03f7a104";
		wait for Clk_period;
		Addr <=  "00001001100111";
		Trees_din <= x"ff7309e5";
		wait for Clk_period;
		Addr <=  "00001001101000";
		Trees_din <= x"06f50204";
		wait for Clk_period;
		Addr <=  "00001001101001";
		Trees_din <= x"ff8109e5";
		wait for Clk_period;
		Addr <=  "00001001101010";
		Trees_din <= x"12febb10";
		wait for Clk_period;
		Addr <=  "00001001101011";
		Trees_din <= x"05feea08";
		wait for Clk_period;
		Addr <=  "00001001101100";
		Trees_din <= x"06f53904";
		wait for Clk_period;
		Addr <=  "00001001101101";
		Trees_din <= x"007309e5";
		wait for Clk_period;
		Addr <=  "00001001101110";
		Trees_din <= x"ffab09e5";
		wait for Clk_period;
		Addr <=  "00001001101111";
		Trees_din <= x"1004d904";
		wait for Clk_period;
		Addr <=  "00001001110000";
		Trees_din <= x"00bd09e5";
		wait for Clk_period;
		Addr <=  "00001001110001";
		Trees_din <= x"000a09e5";
		wait for Clk_period;
		Addr <=  "00001001110010";
		Trees_din <= x"01038908";
		wait for Clk_period;
		Addr <=  "00001001110011";
		Trees_din <= x"0b042604";
		wait for Clk_period;
		Addr <=  "00001001110100";
		Trees_din <= x"000709e5";
		wait for Clk_period;
		Addr <=  "00001001110101";
		Trees_din <= x"ff9c09e5";
		wait for Clk_period;
		Addr <=  "00001001110110";
		Trees_din <= x"07005504";
		wait for Clk_period;
		Addr <=  "00001001110111";
		Trees_din <= x"ffd609e5";
		wait for Clk_period;
		Addr <=  "00001001111000";
		Trees_din <= x"00be09e5";
		wait for Clk_period;
		Addr <=  "00001001111001";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00001001111010";
		Trees_din <= x"05fd340c";
		wait for Clk_period;
		Addr <=  "00001001111011";
		Trees_din <= x"02fc0c08";
		wait for Clk_period;
		Addr <=  "00001001111100";
		Trees_din <= x"10fbfc04";
		wait for Clk_period;
		Addr <=  "00001001111101";
		Trees_din <= x"00450a45";
		wait for Clk_period;
		Addr <=  "00001001111110";
		Trees_din <= x"ffad0a45";
		wait for Clk_period;
		Addr <=  "00001001111111";
		Trees_din <= x"ff680a45";
		wait for Clk_period;
		Addr <=  "00001010000000";
		Trees_din <= x"03f7a104";
		wait for Clk_period;
		Addr <=  "00001010000001";
		Trees_din <= x"ff770a45";
		wait for Clk_period;
		Addr <=  "00001010000010";
		Trees_din <= x"06f50204";
		wait for Clk_period;
		Addr <=  "00001010000011";
		Trees_din <= x"ff850a45";
		wait for Clk_period;
		Addr <=  "00001010000100";
		Trees_din <= x"03f9110c";
		wait for Clk_period;
		Addr <=  "00001010000101";
		Trees_din <= x"0d026504";
		wait for Clk_period;
		Addr <=  "00001010000110";
		Trees_din <= x"ffc60a45";
		wait for Clk_period;
		Addr <=  "00001010000111";
		Trees_din <= x"1700de04";
		wait for Clk_period;
		Addr <=  "00001010001000";
		Trees_din <= x"00180a45";
		wait for Clk_period;
		Addr <=  "00001010001001";
		Trees_din <= x"01350a45";
		wait for Clk_period;
		Addr <=  "00001010001010";
		Trees_din <= x"11fe6008";
		wait for Clk_period;
		Addr <=  "00001010001011";
		Trees_din <= x"0c021b04";
		wait for Clk_period;
		Addr <=  "00001010001100";
		Trees_din <= x"008c0a45";
		wait for Clk_period;
		Addr <=  "00001010001101";
		Trees_din <= x"fff10a45";
		wait for Clk_period;
		Addr <=  "00001010001110";
		Trees_din <= x"0501a404";
		wait for Clk_period;
		Addr <=  "00001010001111";
		Trees_din <= x"ffe50a45";
		wait for Clk_period;
		Addr <=  "00001010010000";
		Trees_din <= x"003d0a45";
		wait for Clk_period;
		Addr <=  "00001010010001";
		Trees_din <= x"05fd4e0c";
		wait for Clk_period;
		Addr <=  "00001010010010";
		Trees_din <= x"07004a04";
		wait for Clk_period;
		Addr <=  "00001010010011";
		Trees_din <= x"fffe0ab1";
		wait for Clk_period;
		Addr <=  "00001010010100";
		Trees_din <= x"05fd3404";
		wait for Clk_period;
		Addr <=  "00001010010101";
		Trees_din <= x"ff690ab1";
		wait for Clk_period;
		Addr <=  "00001010010110";
		Trees_din <= x"ffd00ab1";
		wait for Clk_period;
		Addr <=  "00001010010111";
		Trees_din <= x"03f7a104";
		wait for Clk_period;
		Addr <=  "00001010011000";
		Trees_din <= x"ff7c0ab1";
		wait for Clk_period;
		Addr <=  "00001010011001";
		Trees_din <= x"05040a20";
		wait for Clk_period;
		Addr <=  "00001010011010";
		Trees_din <= x"0e025f10";
		wait for Clk_period;
		Addr <=  "00001010011011";
		Trees_din <= x"05fede08";
		wait for Clk_period;
		Addr <=  "00001010011100";
		Trees_din <= x"00fda604";
		wait for Clk_period;
		Addr <=  "00001010011101";
		Trees_din <= x"001c0ab1";
		wait for Clk_period;
		Addr <=  "00001010011110";
		Trees_din <= x"ff870ab1";
		wait for Clk_period;
		Addr <=  "00001010011111";
		Trees_din <= x"0c024e04";
		wait for Clk_period;
		Addr <=  "00001010100000";
		Trees_din <= x"002b0ab1";
		wait for Clk_period;
		Addr <=  "00001010100001";
		Trees_din <= x"ffb80ab1";
		wait for Clk_period;
		Addr <=  "00001010100010";
		Trees_din <= x"1b003c08";
		wait for Clk_period;
		Addr <=  "00001010100011";
		Trees_din <= x"1d003d04";
		wait for Clk_period;
		Addr <=  "00001010100100";
		Trees_din <= x"ffd50ab1";
		wait for Clk_period;
		Addr <=  "00001010100101";
		Trees_din <= x"009b0ab1";
		wait for Clk_period;
		Addr <=  "00001010100110";
		Trees_din <= x"03fd0604";
		wait for Clk_period;
		Addr <=  "00001010100111";
		Trees_din <= x"ffe00ab1";
		wait for Clk_period;
		Addr <=  "00001010101000";
		Trees_din <= x"ff8a0ab1";
		wait for Clk_period;
		Addr <=  "00001010101001";
		Trees_din <= x"11031f04";
		wait for Clk_period;
		Addr <=  "00001010101010";
		Trees_din <= x"00900ab1";
		wait for Clk_period;
		Addr <=  "00001010101011";
		Trees_din <= x"ffbb0ab1";
		wait for Clk_period;
		Addr <=  "00001010101100";
		Trees_din <= x"05fd3408";
		wait for Clk_period;
		Addr <=  "00001010101101";
		Trees_din <= x"1104aa04";
		wait for Clk_period;
		Addr <=  "00001010101110";
		Trees_din <= x"ff6a0b15";
		wait for Clk_period;
		Addr <=  "00001010101111";
		Trees_din <= x"00080b15";
		wait for Clk_period;
		Addr <=  "00001010110000";
		Trees_din <= x"000fd324";
		wait for Clk_period;
		Addr <=  "00001010110001";
		Trees_din <= x"06f50204";
		wait for Clk_period;
		Addr <=  "00001010110010";
		Trees_din <= x"ff880b15";
		wait for Clk_period;
		Addr <=  "00001010110011";
		Trees_din <= x"01038910";
		wait for Clk_period;
		Addr <=  "00001010110100";
		Trees_din <= x"05fe8a08";
		wait for Clk_period;
		Addr <=  "00001010110101";
		Trees_din <= x"06f76004";
		wait for Clk_period;
		Addr <=  "00001010110110";
		Trees_din <= x"fff70b15";
		wait for Clk_period;
		Addr <=  "00001010110111";
		Trees_din <= x"ff790b15";
		wait for Clk_period;
		Addr <=  "00001010111000";
		Trees_din <= x"11fea804";
		wait for Clk_period;
		Addr <=  "00001010111001";
		Trees_din <= x"00720b15";
		wait for Clk_period;
		Addr <=  "00001010111010";
		Trees_din <= x"00060b15";
		wait for Clk_period;
		Addr <=  "00001010111011";
		Trees_din <= x"1004bf08";
		wait for Clk_period;
		Addr <=  "00001010111100";
		Trees_din <= x"07005504";
		wait for Clk_period;
		Addr <=  "00001010111101";
		Trees_din <= x"ffe80b15";
		wait for Clk_period;
		Addr <=  "00001010111110";
		Trees_din <= x"00ba0b15";
		wait for Clk_period;
		Addr <=  "00001010111111";
		Trees_din <= x"08027004";
		wait for Clk_period;
		Addr <=  "00001011000000";
		Trees_din <= x"ff920b15";
		wait for Clk_period;
		Addr <=  "00001011000001";
		Trees_din <= x"00460b15";
		wait for Clk_period;
		Addr <=  "00001011000010";
		Trees_din <= x"08001004";
		wait for Clk_period;
		Addr <=  "00001011000011";
		Trees_din <= x"00410b15";
		wait for Clk_period;
		Addr <=  "00001011000100";
		Trees_din <= x"ff790b15";
		wait for Clk_period;
		Addr <=  "00001011000101";
		Trees_din <= x"05fd3408";
		wait for Clk_period;
		Addr <=  "00001011000110";
		Trees_din <= x"02fc0c04";
		wait for Clk_period;
		Addr <=  "00001011000111";
		Trees_din <= x"00150b79";
		wait for Clk_period;
		Addr <=  "00001011001000";
		Trees_din <= x"ff6b0b79";
		wait for Clk_period;
		Addr <=  "00001011001001";
		Trees_din <= x"03f7a104";
		wait for Clk_period;
		Addr <=  "00001011001010";
		Trees_din <= x"ff840b79";
		wait for Clk_period;
		Addr <=  "00001011001011";
		Trees_din <= x"03f9110c";
		wait for Clk_period;
		Addr <=  "00001011001100";
		Trees_din <= x"0d026504";
		wait for Clk_period;
		Addr <=  "00001011001101";
		Trees_din <= x"ffc90b79";
		wait for Clk_period;
		Addr <=  "00001011001110";
		Trees_din <= x"1700de04";
		wait for Clk_period;
		Addr <=  "00001011001111";
		Trees_din <= x"00130b79";
		wait for Clk_period;
		Addr <=  "00001011010000";
		Trees_din <= x"00fe0b79";
		wait for Clk_period;
		Addr <=  "00001011010001";
		Trees_din <= x"06f62e0c";
		wait for Clk_period;
		Addr <=  "00001011010010";
		Trees_din <= x"13f8ad04";
		wait for Clk_period;
		Addr <=  "00001011010011";
		Trees_din <= x"00560b79";
		wait for Clk_period;
		Addr <=  "00001011010100";
		Trees_din <= x"05fd5504";
		wait for Clk_period;
		Addr <=  "00001011010101";
		Trees_din <= x"002c0b79";
		wait for Clk_period;
		Addr <=  "00001011010110";
		Trees_din <= x"ff7c0b79";
		wait for Clk_period;
		Addr <=  "00001011010111";
		Trees_din <= x"04fa1608";
		wait for Clk_period;
		Addr <=  "00001011011000";
		Trees_din <= x"0501f804";
		wait for Clk_period;
		Addr <=  "00001011011001";
		Trees_din <= x"ff870b79";
		wait for Clk_period;
		Addr <=  "00001011011010";
		Trees_din <= x"fff70b79";
		wait for Clk_period;
		Addr <=  "00001011011011";
		Trees_din <= x"0e021004";
		wait for Clk_period;
		Addr <=  "00001011011100";
		Trees_din <= x"00000b79";
		wait for Clk_period;
		Addr <=  "00001011011101";
		Trees_din <= x"00480b79";
		wait for Clk_period;
		Addr <=  "00001011011110";
		Trees_din <= x"05fc9304";
		wait for Clk_period;
		Addr <=  "00001011011111";
		Trees_din <= x"ff6c0bd5";
		wait for Clk_period;
		Addr <=  "00001011100000";
		Trees_din <= x"000fd324";
		wait for Clk_period;
		Addr <=  "00001011100001";
		Trees_din <= x"06f50204";
		wait for Clk_period;
		Addr <=  "00001011100010";
		Trees_din <= x"ff8b0bd5";
		wait for Clk_period;
		Addr <=  "00001011100011";
		Trees_din <= x"01038910";
		wait for Clk_period;
		Addr <=  "00001011100100";
		Trees_din <= x"05fe8a08";
		wait for Clk_period;
		Addr <=  "00001011100101";
		Trees_din <= x"09005104";
		wait for Clk_period;
		Addr <=  "00001011100110";
		Trees_din <= x"00070bd5";
		wait for Clk_period;
		Addr <=  "00001011100111";
		Trees_din <= x"ff8e0bd5";
		wait for Clk_period;
		Addr <=  "00001011101000";
		Trees_din <= x"10f8a604";
		wait for Clk_period;
		Addr <=  "00001011101001";
		Trees_din <= x"ffa10bd5";
		wait for Clk_period;
		Addr <=  "00001011101010";
		Trees_din <= x"001f0bd5";
		wait for Clk_period;
		Addr <=  "00001011101011";
		Trees_din <= x"1004bf08";
		wait for Clk_period;
		Addr <=  "00001011101100";
		Trees_din <= x"0bfa0b04";
		wait for Clk_period;
		Addr <=  "00001011101101";
		Trees_din <= x"00fb0bd5";
		wait for Clk_period;
		Addr <=  "00001011101110";
		Trees_din <= x"003f0bd5";
		wait for Clk_period;
		Addr <=  "00001011101111";
		Trees_din <= x"08027004";
		wait for Clk_period;
		Addr <=  "00001011110000";
		Trees_din <= x"ff950bd5";
		wait for Clk_period;
		Addr <=  "00001011110001";
		Trees_din <= x"00400bd5";
		wait for Clk_period;
		Addr <=  "00001011110010";
		Trees_din <= x"06fa7704";
		wait for Clk_period;
		Addr <=  "00001011110011";
		Trees_din <= x"ff7c0bd5";
		wait for Clk_period;
		Addr <=  "00001011110100";
		Trees_din <= x"003d0bd5";
		wait for Clk_period;
		Addr <=  "00001011110101";
		Trees_din <= x"05fc9304";
		wait for Clk_period;
		Addr <=  "00001011110110";
		Trees_din <= x"ff6d0c31";
		wait for Clk_period;
		Addr <=  "00001011110111";
		Trees_din <= x"03f7a104";
		wait for Clk_period;
		Addr <=  "00001011111000";
		Trees_din <= x"ff880c31";
		wait for Clk_period;
		Addr <=  "00001011111001";
		Trees_din <= x"05040a20";
		wait for Clk_period;
		Addr <=  "00001011111010";
		Trees_din <= x"02037010";
		wait for Clk_period;
		Addr <=  "00001011111011";
		Trees_din <= x"08021908";
		wait for Clk_period;
		Addr <=  "00001011111100";
		Trees_din <= x"18004b04";
		wait for Clk_period;
		Addr <=  "00001011111101";
		Trees_din <= x"003c0c31";
		wait for Clk_period;
		Addr <=  "00001011111110";
		Trees_din <= x"ffbc0c31";
		wait for Clk_period;
		Addr <=  "00001011111111";
		Trees_din <= x"18004904";
		wait for Clk_period;
		Addr <=  "00001100000000";
		Trees_din <= x"ffa30c31";
		wait for Clk_period;
		Addr <=  "00001100000001";
		Trees_din <= x"004a0c31";
		wait for Clk_period;
		Addr <=  "00001100000010";
		Trees_din <= x"1b002d08";
		wait for Clk_period;
		Addr <=  "00001100000011";
		Trees_din <= x"1c002904";
		wait for Clk_period;
		Addr <=  "00001100000100";
		Trees_din <= x"00080c31";
		wait for Clk_period;
		Addr <=  "00001100000101";
		Trees_din <= x"00720c31";
		wait for Clk_period;
		Addr <=  "00001100000110";
		Trees_din <= x"09005704";
		wait for Clk_period;
		Addr <=  "00001100000111";
		Trees_din <= x"ff7c0c31";
		wait for Clk_period;
		Addr <=  "00001100001000";
		Trees_din <= x"00060c31";
		wait for Clk_period;
		Addr <=  "00001100001001";
		Trees_din <= x"11031f04";
		wait for Clk_period;
		Addr <=  "00001100001010";
		Trees_din <= x"00860c31";
		wait for Clk_period;
		Addr <=  "00001100001011";
		Trees_din <= x"ffbe0c31";
		wait for Clk_period;
		Addr <=  "00001100001100";
		Trees_din <= x"05fc9304";
		wait for Clk_period;
		Addr <=  "00001100001101";
		Trees_din <= x"ff6f0c8d";
		wait for Clk_period;
		Addr <=  "00001100001110";
		Trees_din <= x"06f50204";
		wait for Clk_period;
		Addr <=  "00001100001111";
		Trees_din <= x"ff8c0c8d";
		wait for Clk_period;
		Addr <=  "00001100010000";
		Trees_din <= x"04f9df0c";
		wait for Clk_period;
		Addr <=  "00001100010001";
		Trees_din <= x"1d005308";
		wait for Clk_period;
		Addr <=  "00001100010010";
		Trees_din <= x"1b003304";
		wait for Clk_period;
		Addr <=  "00001100010011";
		Trees_din <= x"fff20c8d";
		wait for Clk_period;
		Addr <=  "00001100010100";
		Trees_din <= x"ff800c8d";
		wait for Clk_period;
		Addr <=  "00001100010101";
		Trees_din <= x"00450c8d";
		wait for Clk_period;
		Addr <=  "00001100010110";
		Trees_din <= x"11fd5b0c";
		wait for Clk_period;
		Addr <=  "00001100010111";
		Trees_din <= x"18004304";
		wait for Clk_period;
		Addr <=  "00001100011000";
		Trees_din <= x"00010c8d";
		wait for Clk_period;
		Addr <=  "00001100011001";
		Trees_din <= x"09005704";
		wait for Clk_period;
		Addr <=  "00001100011010";
		Trees_din <= x"00ab0c8d";
		wait for Clk_period;
		Addr <=  "00001100011011";
		Trees_din <= x"00210c8d";
		wait for Clk_period;
		Addr <=  "00001100011100";
		Trees_din <= x"0e025f08";
		wait for Clk_period;
		Addr <=  "00001100011101";
		Trees_din <= x"05fede04";
		wait for Clk_period;
		Addr <=  "00001100011110";
		Trees_din <= x"ffaa0c8d";
		wait for Clk_period;
		Addr <=  "00001100011111";
		Trees_din <= x"000e0c8d";
		wait for Clk_period;
		Addr <=  "00001100100000";
		Trees_din <= x"08008504";
		wait for Clk_period;
		Addr <=  "00001100100001";
		Trees_din <= x"ff9c0c8d";
		wait for Clk_period;
		Addr <=  "00001100100010";
		Trees_din <= x"005c0c8d";
		wait for Clk_period;
		Addr <=  "00001100100011";
		Trees_din <= x"05fc9304";
		wait for Clk_period;
		Addr <=  "00001100100100";
		Trees_din <= x"ff700cd9";
		wait for Clk_period;
		Addr <=  "00001100100101";
		Trees_din <= x"06f50204";
		wait for Clk_period;
		Addr <=  "00001100100110";
		Trees_din <= x"ff900cd9";
		wait for Clk_period;
		Addr <=  "00001100100111";
		Trees_din <= x"000fd318";
		wait for Clk_period;
		Addr <=  "00001100101000";
		Trees_din <= x"11fd5b08";
		wait for Clk_period;
		Addr <=  "00001100101001";
		Trees_din <= x"18004304";
		wait for Clk_period;
		Addr <=  "00001100101010";
		Trees_din <= x"00080cd9";
		wait for Clk_period;
		Addr <=  "00001100101011";
		Trees_din <= x"008c0cd9";
		wait for Clk_period;
		Addr <=  "00001100101100";
		Trees_din <= x"01041b08";
		wait for Clk_period;
		Addr <=  "00001100101101";
		Trees_din <= x"0500f004";
		wait for Clk_period;
		Addr <=  "00001100101110";
		Trees_din <= x"ffd60cd9";
		wait for Clk_period;
		Addr <=  "00001100101111";
		Trees_din <= x"002d0cd9";
		wait for Clk_period;
		Addr <=  "00001100110000";
		Trees_din <= x"08009104";
		wait for Clk_period;
		Addr <=  "00001100110001";
		Trees_din <= x"ffd30cd9";
		wait for Clk_period;
		Addr <=  "00001100110010";
		Trees_din <= x"00780cd9";
		wait for Clk_period;
		Addr <=  "00001100110011";
		Trees_din <= x"09004c04";
		wait for Clk_period;
		Addr <=  "00001100110100";
		Trees_din <= x"003c0cd9";
		wait for Clk_period;
		Addr <=  "00001100110101";
		Trees_din <= x"ff870cd9";
		wait for Clk_period;
		Addr <=  "00001100110110";
		Trees_din <= x"05fc9304";
		wait for Clk_period;
		Addr <=  "00001100110111";
		Trees_din <= x"ff720d85";
		wait for Clk_period;
		Addr <=  "00001100111000";
		Trees_din <= x"0700572c";
		wait for Clk_period;
		Addr <=  "00001100111001";
		Trees_din <= x"0d03171c";
		wait for Clk_period;
		Addr <=  "00001100111010";
		Trees_din <= x"11fe960c";
		wait for Clk_period;
		Addr <=  "00001100111011";
		Trees_din <= x"1e006708";
		wait for Clk_period;
		Addr <=  "00001100111100";
		Trees_din <= x"02014b04";
		wait for Clk_period;
		Addr <=  "00001100111101";
		Trees_din <= x"fffe0d85";
		wait for Clk_period;
		Addr <=  "00001100111110";
		Trees_din <= x"00120d85";
		wait for Clk_period;
		Addr <=  "00001100111111";
		Trees_din <= x"00810d85";
		wait for Clk_period;
		Addr <=  "00001101000000";
		Trees_din <= x"0c02f908";
		wait for Clk_period;
		Addr <=  "00001101000001";
		Trees_din <= x"07005604";
		wait for Clk_period;
		Addr <=  "00001101000010";
		Trees_din <= x"ffba0d85";
		wait for Clk_period;
		Addr <=  "00001101000011";
		Trees_din <= x"002b0d85";
		wait for Clk_period;
		Addr <=  "00001101000100";
		Trees_din <= x"07004a04";
		wait for Clk_period;
		Addr <=  "00001101000101";
		Trees_din <= x"00a60d85";
		wait for Clk_period;
		Addr <=  "00001101000110";
		Trees_din <= x"fffa0d85";
		wait for Clk_period;
		Addr <=  "00001101000111";
		Trees_din <= x"17003204";
		wait for Clk_period;
		Addr <=  "00001101001000";
		Trees_din <= x"ffab0d85";
		wait for Clk_period;
		Addr <=  "00001101001001";
		Trees_din <= x"1500a408";
		wait for Clk_period;
		Addr <=  "00001101001010";
		Trees_din <= x"1a00c104";
		wait for Clk_period;
		Addr <=  "00001101001011";
		Trees_din <= x"00310d85";
		wait for Clk_period;
		Addr <=  "00001101001100";
		Trees_din <= x"00ba0d85";
		wait for Clk_period;
		Addr <=  "00001101001101";
		Trees_din <= x"ffe70d85";
		wait for Clk_period;
		Addr <=  "00001101001110";
		Trees_din <= x"1301ab20";
		wait for Clk_period;
		Addr <=  "00001101001111";
		Trees_din <= x"17031510";
		wait for Clk_period;
		Addr <=  "00001101010000";
		Trees_din <= x"05024c08";
		wait for Clk_period;
		Addr <=  "00001101010001";
		Trees_din <= x"0c037804";
		wait for Clk_period;
		Addr <=  "00001101010010";
		Trees_din <= x"ff7f0d85";
		wait for Clk_period;
		Addr <=  "00001101010011";
		Trees_din <= x"000d0d85";
		wait for Clk_period;
		Addr <=  "00001101010100";
		Trees_din <= x"0e008204";
		wait for Clk_period;
		Addr <=  "00001101010101";
		Trees_din <= x"005f0d85";
		wait for Clk_period;
		Addr <=  "00001101010110";
		Trees_din <= x"ffd80d85";
		wait for Clk_period;
		Addr <=  "00001101010111";
		Trees_din <= x"00feb708";
		wait for Clk_period;
		Addr <=  "00001101011000";
		Trees_din <= x"11012204";
		wait for Clk_period;
		Addr <=  "00001101011001";
		Trees_din <= x"ffff0d85";
		wait for Clk_period;
		Addr <=  "00001101011010";
		Trees_din <= x"008b0d85";
		wait for Clk_period;
		Addr <=  "00001101011011";
		Trees_din <= x"06f83404";
		wait for Clk_period;
		Addr <=  "00001101011100";
		Trees_din <= x"ff9d0d85";
		wait for Clk_period;
		Addr <=  "00001101011101";
		Trees_din <= x"00170d85";
		wait for Clk_period;
		Addr <=  "00001101011110";
		Trees_din <= x"0c010104";
		wait for Clk_period;
		Addr <=  "00001101011111";
		Trees_din <= x"00710d85";
		wait for Clk_period;
		Addr <=  "00001101100000";
		Trees_din <= x"00050d85";
		wait for Clk_period;
		Addr <=  "00001101100001";
		Trees_din <= x"05fc9304";
		wait for Clk_period;
		Addr <=  "00001101100010";
		Trees_din <= x"ff740e31";
		wait for Clk_period;
		Addr <=  "00001101100011";
		Trees_din <= x"0500582c";
		wait for Clk_period;
		Addr <=  "00001101100100";
		Trees_din <= x"02036320";
		wait for Clk_period;
		Addr <=  "00001101100101";
		Trees_din <= x"1e006710";
		wait for Clk_period;
		Addr <=  "00001101100110";
		Trees_din <= x"0afcc208";
		wait for Clk_period;
		Addr <=  "00001101100111";
		Trees_din <= x"17024204";
		wait for Clk_period;
		Addr <=  "00001101101000";
		Trees_din <= x"00500e31";
		wait for Clk_period;
		Addr <=  "00001101101001";
		Trees_din <= x"ffc00e31";
		wait for Clk_period;
		Addr <=  "00001101101010";
		Trees_din <= x"11fd0404";
		wait for Clk_period;
		Addr <=  "00001101101011";
		Trees_din <= x"ffe90e31";
		wait for Clk_period;
		Addr <=  "00001101101100";
		Trees_din <= x"ff730e31";
		wait for Clk_period;
		Addr <=  "00001101101101";
		Trees_din <= x"1a00c808";
		wait for Clk_period;
		Addr <=  "00001101101110";
		Trees_din <= x"15009304";
		wait for Clk_period;
		Addr <=  "00001101101111";
		Trees_din <= x"ffc40e31";
		wait for Clk_period;
		Addr <=  "00001101110000";
		Trees_din <= x"00410e31";
		wait for Clk_period;
		Addr <=  "00001101110001";
		Trees_din <= x"13ff6704";
		wait for Clk_period;
		Addr <=  "00001101110010";
		Trees_din <= x"00170e31";
		wait for Clk_period;
		Addr <=  "00001101110011";
		Trees_din <= x"00c00e31";
		wait for Clk_period;
		Addr <=  "00001101110100";
		Trees_din <= x"01042f04";
		wait for Clk_period;
		Addr <=  "00001101110101";
		Trees_din <= x"ff770e31";
		wait for Clk_period;
		Addr <=  "00001101110110";
		Trees_din <= x"0801d404";
		wait for Clk_period;
		Addr <=  "00001101110111";
		Trees_din <= x"ffab0e31";
		wait for Clk_period;
		Addr <=  "00001101111000";
		Trees_din <= x"00710e31";
		wait for Clk_period;
		Addr <=  "00001101111001";
		Trees_din <= x"13ffb118";
		wait for Clk_period;
		Addr <=  "00001101111010";
		Trees_din <= x"0700590c";
		wait for Clk_period;
		Addr <=  "00001101111011";
		Trees_din <= x"11028708";
		wait for Clk_period;
		Addr <=  "00001101111100";
		Trees_din <= x"01fb5b04";
		wait for Clk_period;
		Addr <=  "00001101111101";
		Trees_din <= x"00050e31";
		wait for Clk_period;
		Addr <=  "00001101111110";
		Trees_din <= x"00860e31";
		wait for Clk_period;
		Addr <=  "00001101111111";
		Trees_din <= x"ffdb0e31";
		wait for Clk_period;
		Addr <=  "00001110000000";
		Trees_din <= x"19008c04";
		wait for Clk_period;
		Addr <=  "00001110000001";
		Trees_din <= x"00470e31";
		wait for Clk_period;
		Addr <=  "00001110000010";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00001110000011";
		Trees_din <= x"ffa10e31";
		wait for Clk_period;
		Addr <=  "00001110000100";
		Trees_din <= x"ffe90e31";
		wait for Clk_period;
		Addr <=  "00001110000101";
		Trees_din <= x"15009e08";
		wait for Clk_period;
		Addr <=  "00001110000110";
		Trees_din <= x"18004804";
		wait for Clk_period;
		Addr <=  "00001110000111";
		Trees_din <= x"ff940e31";
		wait for Clk_period;
		Addr <=  "00001110001000";
		Trees_din <= x"00230e31";
		wait for Clk_period;
		Addr <=  "00001110001001";
		Trees_din <= x"10fba804";
		wait for Clk_period;
		Addr <=  "00001110001010";
		Trees_din <= x"00420e31";
		wait for Clk_period;
		Addr <=  "00001110001011";
		Trees_din <= x"fffa0e31";
		wait for Clk_period;
		Addr <=  "00001110001100";
		Trees_din <= x"05fc9304";
		wait for Clk_period;
		Addr <=  "00001110001101";
		Trees_din <= x"ff760e9d";
		wait for Clk_period;
		Addr <=  "00001110001110";
		Trees_din <= x"06f50204";
		wait for Clk_period;
		Addr <=  "00001110001111";
		Trees_din <= x"ff990e9d";
		wait for Clk_period;
		Addr <=  "00001110010000";
		Trees_din <= x"04fb5414";
		wait for Clk_period;
		Addr <=  "00001110010001";
		Trees_din <= x"0503440c";
		wait for Clk_period;
		Addr <=  "00001110010010";
		Trees_din <= x"1a00b708";
		wait for Clk_period;
		Addr <=  "00001110010011";
		Trees_din <= x"1c003e04";
		wait for Clk_period;
		Addr <=  "00001110010100";
		Trees_din <= x"004c0e9d";
		wait for Clk_period;
		Addr <=  "00001110010101";
		Trees_din <= x"ffc10e9d";
		wait for Clk_period;
		Addr <=  "00001110010110";
		Trees_din <= x"ff7d0e9d";
		wait for Clk_period;
		Addr <=  "00001110010111";
		Trees_din <= x"08008c04";
		wait for Clk_period;
		Addr <=  "00001110011000";
		Trees_din <= x"ffe20e9d";
		wait for Clk_period;
		Addr <=  "00001110011001";
		Trees_din <= x"00520e9d";
		wait for Clk_period;
		Addr <=  "00001110011010";
		Trees_din <= x"1400fa10";
		wait for Clk_period;
		Addr <=  "00001110011011";
		Trees_din <= x"07005808";
		wait for Clk_period;
		Addr <=  "00001110011100";
		Trees_din <= x"17028804";
		wait for Clk_period;
		Addr <=  "00001110011101";
		Trees_din <= x"00720e9d";
		wait for Clk_period;
		Addr <=  "00001110011110";
		Trees_din <= x"00060e9d";
		wait for Clk_period;
		Addr <=  "00001110011111";
		Trees_din <= x"00feb704";
		wait for Clk_period;
		Addr <=  "00001110100000";
		Trees_din <= x"00380e9d";
		wait for Clk_period;
		Addr <=  "00001110100001";
		Trees_din <= x"ffa10e9d";
		wait for Clk_period;
		Addr <=  "00001110100010";
		Trees_din <= x"0305c708";
		wait for Clk_period;
		Addr <=  "00001110100011";
		Trees_din <= x"15009b04";
		wait for Clk_period;
		Addr <=  "00001110100100";
		Trees_din <= x"00330e9d";
		wait for Clk_period;
		Addr <=  "00001110100101";
		Trees_din <= x"ffd10e9d";
		wait for Clk_period;
		Addr <=  "00001110100110";
		Trees_din <= x"ff840e9d";
		wait for Clk_period;
		Addr <=  "00001110100111";
		Trees_din <= x"05fc9304";
		wait for Clk_period;
		Addr <=  "00001110101000";
		Trees_din <= x"ff780f41";
		wait for Clk_period;
		Addr <=  "00001110101001";
		Trees_din <= x"05005834";
		wait for Clk_period;
		Addr <=  "00001110101010";
		Trees_din <= x"0c008c14";
		wait for Clk_period;
		Addr <=  "00001110101011";
		Trees_din <= x"14003308";
		wait for Clk_period;
		Addr <=  "00001110101100";
		Trees_din <= x"11007904";
		wait for Clk_period;
		Addr <=  "00001110101101";
		Trees_din <= x"ffea0f41";
		wait for Clk_period;
		Addr <=  "00001110101110";
		Trees_din <= x"ffa90f41";
		wait for Clk_period;
		Addr <=  "00001110101111";
		Trees_din <= x"1403e008";
		wait for Clk_period;
		Addr <=  "00001110110000";
		Trees_din <= x"13fdaa04";
		wait for Clk_period;
		Addr <=  "00001110110001";
		Trees_din <= x"002a0f41";
		wait for Clk_period;
		Addr <=  "00001110110010";
		Trees_din <= x"009b0f41";
		wait for Clk_period;
		Addr <=  "00001110110011";
		Trees_din <= x"ffc10f41";
		wait for Clk_period;
		Addr <=  "00001110110100";
		Trees_din <= x"02ffbf10";
		wait for Clk_period;
		Addr <=  "00001110110101";
		Trees_din <= x"0b027508";
		wait for Clk_period;
		Addr <=  "00001110110110";
		Trees_din <= x"1a00c204";
		wait for Clk_period;
		Addr <=  "00001110110111";
		Trees_din <= x"ffa70f41";
		wait for Clk_period;
		Addr <=  "00001110111000";
		Trees_din <= x"006e0f41";
		wait for Clk_period;
		Addr <=  "00001110111001";
		Trees_din <= x"08009104";
		wait for Clk_period;
		Addr <=  "00001110111010";
		Trees_din <= x"00240f41";
		wait for Clk_period;
		Addr <=  "00001110111011";
		Trees_din <= x"ff800f41";
		wait for Clk_period;
		Addr <=  "00001110111100";
		Trees_din <= x"11fe6008";
		wait for Clk_period;
		Addr <=  "00001110111101";
		Trees_din <= x"19008e04";
		wait for Clk_period;
		Addr <=  "00001110111110";
		Trees_din <= x"005b0f41";
		wait for Clk_period;
		Addr <=  "00001110111111";
		Trees_din <= x"ffd60f41";
		wait for Clk_period;
		Addr <=  "00001111000000";
		Trees_din <= x"06f82604";
		wait for Clk_period;
		Addr <=  "00001111000001";
		Trees_din <= x"ff6f0f41";
		wait for Clk_period;
		Addr <=  "00001111000010";
		Trees_din <= x"ffe30f41";
		wait for Clk_period;
		Addr <=  "00001111000011";
		Trees_din <= x"12028714";
		wait for Clk_period;
		Addr <=  "00001111000100";
		Trees_din <= x"1004ce0c";
		wait for Clk_period;
		Addr <=  "00001111000101";
		Trees_din <= x"10f92b04";
		wait for Clk_period;
		Addr <=  "00001111000110";
		Trees_din <= x"ffdd0f41";
		wait for Clk_period;
		Addr <=  "00001111000111";
		Trees_din <= x"0801ca04";
		wait for Clk_period;
		Addr <=  "00001111001000";
		Trees_din <= x"007d0f41";
		wait for Clk_period;
		Addr <=  "00001111001001";
		Trees_din <= x"001d0f41";
		wait for Clk_period;
		Addr <=  "00001111001010";
		Trees_din <= x"0f016804";
		wait for Clk_period;
		Addr <=  "00001111001011";
		Trees_din <= x"ffa00f41";
		wait for Clk_period;
		Addr <=  "00001111001100";
		Trees_din <= x"00420f41";
		wait for Clk_period;
		Addr <=  "00001111001101";
		Trees_din <= x"19009504";
		wait for Clk_period;
		Addr <=  "00001111001110";
		Trees_din <= x"ffa70f41";
		wait for Clk_period;
		Addr <=  "00001111001111";
		Trees_din <= x"00240f41";
		wait for Clk_period;
		Addr <=  "00001111010000";
		Trees_din <= x"05fc9304";
		wait for Clk_period;
		Addr <=  "00001111010001";
		Trees_din <= x"ff7b0fed";
		wait for Clk_period;
		Addr <=  "00001111010010";
		Trees_din <= x"00068130";
		wait for Clk_period;
		Addr <=  "00001111010011";
		Trees_din <= x"01fec714";
		wait for Clk_period;
		Addr <=  "00001111010100";
		Trees_din <= x"0900580c";
		wait for Clk_period;
		Addr <=  "00001111010101";
		Trees_din <= x"1c002a04";
		wait for Clk_period;
		Addr <=  "00001111010110";
		Trees_din <= x"ff9e0fed";
		wait for Clk_period;
		Addr <=  "00001111010111";
		Trees_din <= x"1401a404";
		wait for Clk_period;
		Addr <=  "00001111011000";
		Trees_din <= x"00590fed";
		wait for Clk_period;
		Addr <=  "00001111011001";
		Trees_din <= x"fff40fed";
		wait for Clk_period;
		Addr <=  "00001111011010";
		Trees_din <= x"0d030d04";
		wait for Clk_period;
		Addr <=  "00001111011011";
		Trees_din <= x"ff8b0fed";
		wait for Clk_period;
		Addr <=  "00001111011100";
		Trees_din <= x"ffff0fed";
		wait for Clk_period;
		Addr <=  "00001111011101";
		Trees_din <= x"05feea0c";
		wait for Clk_period;
		Addr <=  "00001111011110";
		Trees_din <= x"01038904";
		wait for Clk_period;
		Addr <=  "00001111011111";
		Trees_din <= x"ff910fed";
		wait for Clk_period;
		Addr <=  "00001111100000";
		Trees_din <= x"03fe8b04";
		wait for Clk_period;
		Addr <=  "00001111100001";
		Trees_din <= x"ffc50fed";
		wait for Clk_period;
		Addr <=  "00001111100010";
		Trees_din <= x"00660fed";
		wait for Clk_period;
		Addr <=  "00001111100011";
		Trees_din <= x"06f66908";
		wait for Clk_period;
		Addr <=  "00001111100100";
		Trees_din <= x"0b04c704";
		wait for Clk_period;
		Addr <=  "00001111100101";
		Trees_din <= x"ffcd0fed";
		wait for Clk_period;
		Addr <=  "00001111100110";
		Trees_din <= x"00550fed";
		wait for Clk_period;
		Addr <=  "00001111100111";
		Trees_din <= x"0f001904";
		wait for Clk_period;
		Addr <=  "00001111101000";
		Trees_din <= x"000b0fed";
		wait for Clk_period;
		Addr <=  "00001111101001";
		Trees_din <= x"00870fed";
		wait for Clk_period;
		Addr <=  "00001111101010";
		Trees_din <= x"0a038918";
		wait for Clk_period;
		Addr <=  "00001111101011";
		Trees_din <= x"0500f008";
		wait for Clk_period;
		Addr <=  "00001111101100";
		Trees_din <= x"1403c904";
		wait for Clk_period;
		Addr <=  "00001111101101";
		Trees_din <= x"ff780fed";
		wait for Clk_period;
		Addr <=  "00001111101110";
		Trees_din <= x"001c0fed";
		wait for Clk_period;
		Addr <=  "00001111101111";
		Trees_din <= x"13fe5a08";
		wait for Clk_period;
		Addr <=  "00001111110000";
		Trees_din <= x"16038f04";
		wait for Clk_period;
		Addr <=  "00001111110001";
		Trees_din <= x"00180fed";
		wait for Clk_period;
		Addr <=  "00001111110010";
		Trees_din <= x"00510fed";
		wait for Clk_period;
		Addr <=  "00001111110011";
		Trees_din <= x"09005604";
		wait for Clk_period;
		Addr <=  "00001111110100";
		Trees_din <= x"ffac0fed";
		wait for Clk_period;
		Addr <=  "00001111110101";
		Trees_din <= x"00260fed";
		wait for Clk_period;
		Addr <=  "00001111110110";
		Trees_din <= x"0a03b704";
		wait for Clk_period;
		Addr <=  "00001111110111";
		Trees_din <= x"00920fed";
		wait for Clk_period;
		Addr <=  "00001111111000";
		Trees_din <= x"0009f004";
		wait for Clk_period;
		Addr <=  "00001111111001";
		Trees_din <= x"000f0fed";
		wait for Clk_period;
		Addr <=  "00001111111010";
		Trees_din <= x"ffad0fed";
		wait for Clk_period;
		Addr <=  "00001111111011";
		Trees_din <= x"05fc9304";
		wait for Clk_period;
		Addr <=  "00001111111100";
		Trees_din <= x"ff7e1069";
		wait for Clk_period;
		Addr <=  "00001111111101";
		Trees_din <= x"12febb18";
		wait for Clk_period;
		Addr <=  "00001111111110";
		Trees_din <= x"05feea08";
		wait for Clk_period;
		Addr <=  "00001111111111";
		Trees_din <= x"13fe5104";
		wait for Clk_period;
		Addr <=  "00010000000000";
		Trees_din <= x"ffad1069";
		wait for Clk_period;
		Addr <=  "00010000000001";
		Trees_din <= x"001a1069";
		wait for Clk_period;
		Addr <=  "00010000000010";
		Trees_din <= x"1004d908";
		wait for Clk_period;
		Addr <=  "00010000000011";
		Trees_din <= x"01001f04";
		wait for Clk_period;
		Addr <=  "00010000000100";
		Trees_din <= x"00851069";
		wait for Clk_period;
		Addr <=  "00010000000101";
		Trees_din <= x"001a1069";
		wait for Clk_period;
		Addr <=  "00010000000110";
		Trees_din <= x"01fd2104";
		wait for Clk_period;
		Addr <=  "00010000000111";
		Trees_din <= x"00351069";
		wait for Clk_period;
		Addr <=  "00010000001000";
		Trees_din <= x"ffb61069";
		wait for Clk_period;
		Addr <=  "00010000001001";
		Trees_din <= x"12003308";
		wait for Clk_period;
		Addr <=  "00010000001010";
		Trees_din <= x"04fcef04";
		wait for Clk_period;
		Addr <=  "00010000001011";
		Trees_din <= x"ffea1069";
		wait for Clk_period;
		Addr <=  "00010000001100";
		Trees_din <= x"ff861069";
		wait for Clk_period;
		Addr <=  "00010000001101";
		Trees_din <= x"1a00c20c";
		wait for Clk_period;
		Addr <=  "00010000001110";
		Trees_din <= x"0c024108";
		wait for Clk_period;
		Addr <=  "00010000001111";
		Trees_din <= x"05007904";
		wait for Clk_period;
		Addr <=  "00010000010000";
		Trees_din <= x"ffd11069";
		wait for Clk_period;
		Addr <=  "00010000010001";
		Trees_din <= x"00311069";
		wait for Clk_period;
		Addr <=  "00010000010010";
		Trees_din <= x"ff851069";
		wait for Clk_period;
		Addr <=  "00010000010011";
		Trees_din <= x"1c003308";
		wait for Clk_period;
		Addr <=  "00010000010100";
		Trees_din <= x"05009b04";
		wait for Clk_period;
		Addr <=  "00010000010101";
		Trees_din <= x"ffcc1069";
		wait for Clk_period;
		Addr <=  "00010000010110";
		Trees_din <= x"00221069";
		wait for Clk_period;
		Addr <=  "00010000010111";
		Trees_din <= x"04fe1204";
		wait for Clk_period;
		Addr <=  "00010000011000";
		Trees_din <= x"ffaf1069";
		wait for Clk_period;
		Addr <=  "00010000011001";
		Trees_din <= x"00861069";
		wait for Clk_period;
		Addr <=  "00010000011010";
		Trees_din <= x"05fc9304";
		wait for Clk_period;
		Addr <=  "00010000011011";
		Trees_din <= x"ff8010c5";
		wait for Clk_period;
		Addr <=  "00010000011100";
		Trees_din <= x"05040a24";
		wait for Clk_period;
		Addr <=  "00010000011101";
		Trees_din <= x"02037010";
		wait for Clk_period;
		Addr <=  "00010000011110";
		Trees_din <= x"0efbda04";
		wait for Clk_period;
		Addr <=  "00010000011111";
		Trees_din <= x"ffaa10c5";
		wait for Clk_period;
		Addr <=  "00010000100000";
		Trees_din <= x"04fac204";
		wait for Clk_period;
		Addr <=  "00010000100001";
		Trees_din <= x"ffad10c5";
		wait for Clk_period;
		Addr <=  "00010000100010";
		Trees_din <= x"1a00f404";
		wait for Clk_period;
		Addr <=  "00010000100011";
		Trees_din <= x"002c10c5";
		wait for Clk_period;
		Addr <=  "00010000100100";
		Trees_din <= x"ffc210c5";
		wait for Clk_period;
		Addr <=  "00010000100101";
		Trees_din <= x"1b002d04";
		wait for Clk_period;
		Addr <=  "00010000100110";
		Trees_din <= x"003810c5";
		wait for Clk_period;
		Addr <=  "00010000100111";
		Trees_din <= x"09005708";
		wait for Clk_period;
		Addr <=  "00010000101000";
		Trees_din <= x"17000004";
		wait for Clk_period;
		Addr <=  "00010000101001";
		Trees_din <= x"ffd710c5";
		wait for Clk_period;
		Addr <=  "00010000101010";
		Trees_din <= x"ff7b10c5";
		wait for Clk_period;
		Addr <=  "00010000101011";
		Trees_din <= x"07005704";
		wait for Clk_period;
		Addr <=  "00010000101100";
		Trees_din <= x"004410c5";
		wait for Clk_period;
		Addr <=  "00010000101101";
		Trees_din <= x"ffc310c5";
		wait for Clk_period;
		Addr <=  "00010000101110";
		Trees_din <= x"0e026504";
		wait for Clk_period;
		Addr <=  "00010000101111";
		Trees_din <= x"005a10c5";
		wait for Clk_period;
		Addr <=  "00010000110000";
		Trees_din <= x"fff310c5";
		wait for Clk_period;
		Addr <=  "00010000110001";
		Trees_din <= x"05fc9304";
		wait for Clk_period;
		Addr <=  "00010000110010";
		Trees_din <= x"ff841131";
		wait for Clk_period;
		Addr <=  "00010000110011";
		Trees_din <= x"1c002208";
		wait for Clk_period;
		Addr <=  "00010000110100";
		Trees_din <= x"0b03ea04";
		wait for Clk_period;
		Addr <=  "00010000110101";
		Trees_din <= x"ffe41131";
		wait for Clk_period;
		Addr <=  "00010000110110";
		Trees_din <= x"007b1131";
		wait for Clk_period;
		Addr <=  "00010000110111";
		Trees_din <= x"1c002d10";
		wait for Clk_period;
		Addr <=  "00010000111000";
		Trees_din <= x"1b002c08";
		wait for Clk_period;
		Addr <=  "00010000111001";
		Trees_din <= x"18003504";
		wait for Clk_period;
		Addr <=  "00010000111010";
		Trees_din <= x"ffb01131";
		wait for Clk_period;
		Addr <=  "00010000111011";
		Trees_din <= x"005d1131";
		wait for Clk_period;
		Addr <=  "00010000111100";
		Trees_din <= x"0d00ae04";
		wait for Clk_period;
		Addr <=  "00010000111101";
		Trees_din <= x"ffe11131";
		wait for Clk_period;
		Addr <=  "00010000111110";
		Trees_din <= x"ff811131";
		wait for Clk_period;
		Addr <=  "00010000111111";
		Trees_din <= x"08006810";
		wait for Clk_period;
		Addr <=  "00010001000000";
		Trees_din <= x"1b004508";
		wait for Clk_period;
		Addr <=  "00010001000001";
		Trees_din <= x"1c003204";
		wait for Clk_period;
		Addr <=  "00010001000010";
		Trees_din <= x"00021131";
		wait for Clk_period;
		Addr <=  "00010001000011";
		Trees_din <= x"ff841131";
		wait for Clk_period;
		Addr <=  "00010001000100";
		Trees_din <= x"1200a404";
		wait for Clk_period;
		Addr <=  "00010001000101";
		Trees_din <= x"004a1131";
		wait for Clk_period;
		Addr <=  "00010001000110";
		Trees_din <= x"ffc31131";
		wait for Clk_period;
		Addr <=  "00010001000111";
		Trees_din <= x"08009304";
		wait for Clk_period;
		Addr <=  "00010001001000";
		Trees_din <= x"00731131";
		wait for Clk_period;
		Addr <=  "00010001001001";
		Trees_din <= x"06f66f04";
		wait for Clk_period;
		Addr <=  "00010001001010";
		Trees_din <= x"ffae1131";
		wait for Clk_period;
		Addr <=  "00010001001011";
		Trees_din <= x"001a1131";
		wait for Clk_period;
		Addr <=  "00010001001100";
		Trees_din <= x"05fc9304";
		wait for Clk_period;
		Addr <=  "00010001001101";
		Trees_din <= x"ff8711bd";
		wait for Clk_period;
		Addr <=  "00010001001110";
		Trees_din <= x"00015520";
		wait for Clk_period;
		Addr <=  "00010001001111";
		Trees_din <= x"13ffcc14";
		wait for Clk_period;
		Addr <=  "00010001010000";
		Trees_din <= x"05fe1004";
		wait for Clk_period;
		Addr <=  "00010001010001";
		Trees_din <= x"ff9d11bd";
		wait for Clk_period;
		Addr <=  "00010001010010";
		Trees_din <= x"17027908";
		wait for Clk_period;
		Addr <=  "00010001010011";
		Trees_din <= x"0c02eb04";
		wait for Clk_period;
		Addr <=  "00010001010100";
		Trees_din <= x"ff9311bd";
		wait for Clk_period;
		Addr <=  "00010001010101";
		Trees_din <= x"004e11bd";
		wait for Clk_period;
		Addr <=  "00010001010110";
		Trees_din <= x"1d004304";
		wait for Clk_period;
		Addr <=  "00010001010111";
		Trees_din <= x"001d11bd";
		wait for Clk_period;
		Addr <=  "00010001011000";
		Trees_din <= x"006a11bd";
		wait for Clk_period;
		Addr <=  "00010001011001";
		Trees_din <= x"01fd3904";
		wait for Clk_period;
		Addr <=  "00010001011010";
		Trees_din <= x"ffde11bd";
		wait for Clk_period;
		Addr <=  "00010001011011";
		Trees_din <= x"1c002d04";
		wait for Clk_period;
		Addr <=  "00010001011100";
		Trees_din <= x"000911bd";
		wait for Clk_period;
		Addr <=  "00010001011101";
		Trees_din <= x"008311bd";
		wait for Clk_period;
		Addr <=  "00010001011110";
		Trees_din <= x"12fe9910";
		wait for Clk_period;
		Addr <=  "00010001011111";
		Trees_din <= x"0700570c";
		wait for Clk_period;
		Addr <=  "00010001100000";
		Trees_din <= x"09005508";
		wait for Clk_period;
		Addr <=  "00010001100001";
		Trees_din <= x"06f87f04";
		wait for Clk_period;
		Addr <=  "00010001100010";
		Trees_din <= x"002311bd";
		wait for Clk_period;
		Addr <=  "00010001100011";
		Trees_din <= x"007c11bd";
		wait for Clk_period;
		Addr <=  "00010001100100";
		Trees_din <= x"fff711bd";
		wait for Clk_period;
		Addr <=  "00010001100101";
		Trees_din <= x"ffe011bd";
		wait for Clk_period;
		Addr <=  "00010001100110";
		Trees_din <= x"1200e704";
		wait for Clk_period;
		Addr <=  "00010001100111";
		Trees_din <= x"ff9411bd";
		wait for Clk_period;
		Addr <=  "00010001101000";
		Trees_din <= x"15009508";
		wait for Clk_period;
		Addr <=  "00010001101001";
		Trees_din <= x"0e003904";
		wait for Clk_period;
		Addr <=  "00010001101010";
		Trees_din <= x"001a11bd";
		wait for Clk_period;
		Addr <=  "00010001101011";
		Trees_din <= x"ff9111bd";
		wait for Clk_period;
		Addr <=  "00010001101100";
		Trees_din <= x"1b003304";
		wait for Clk_period;
		Addr <=  "00010001101101";
		Trees_din <= x"ffd711bd";
		wait for Clk_period;
		Addr <=  "00010001101110";
		Trees_din <= x"004c11bd";
		wait for Clk_period;
		Addr <=  "00010001101111";
		Trees_din <= x"05fc9304";
		wait for Clk_period;
		Addr <=  "00010001110000";
		Trees_din <= x"ff8b1259";
		wait for Clk_period;
		Addr <=  "00010001110001";
		Trees_din <= x"05005828";
		wait for Clk_period;
		Addr <=  "00010001110010";
		Trees_din <= x"0c012a14";
		wait for Clk_period;
		Addr <=  "00010001110011";
		Trees_din <= x"13fd8c08";
		wait for Clk_period;
		Addr <=  "00010001110100";
		Trees_din <= x"05feea04";
		wait for Clk_period;
		Addr <=  "00010001110101";
		Trees_din <= x"ff9f1259";
		wait for Clk_period;
		Addr <=  "00010001110110";
		Trees_din <= x"000c1259";
		wait for Clk_period;
		Addr <=  "00010001110111";
		Trees_din <= x"02036308";
		wait for Clk_period;
		Addr <=  "00010001111000";
		Trees_din <= x"18004904";
		wait for Clk_period;
		Addr <=  "00010001111001";
		Trees_din <= x"006a1259";
		wait for Clk_period;
		Addr <=  "00010001111010";
		Trees_din <= x"ffcc1259";
		wait for Clk_period;
		Addr <=  "00010001111011";
		Trees_din <= x"ffb01259";
		wait for Clk_period;
		Addr <=  "00010001111100";
		Trees_din <= x"03029108";
		wait for Clk_period;
		Addr <=  "00010001111101";
		Trees_din <= x"0d00bc04";
		wait for Clk_period;
		Addr <=  "00010001111110";
		Trees_din <= x"fffc1259";
		wait for Clk_period;
		Addr <=  "00010001111111";
		Trees_din <= x"ff851259";
		wait for Clk_period;
		Addr <=  "00010010000000";
		Trees_din <= x"0b027508";
		wait for Clk_period;
		Addr <=  "00010010000001";
		Trees_din <= x"01fd3904";
		wait for Clk_period;
		Addr <=  "00010010000010";
		Trees_din <= x"ffd81259";
		wait for Clk_period;
		Addr <=  "00010010000011";
		Trees_din <= x"00651259";
		wait for Clk_period;
		Addr <=  "00010010000100";
		Trees_din <= x"ffa81259";
		wait for Clk_period;
		Addr <=  "00010010000101";
		Trees_din <= x"06f9ff18";
		wait for Clk_period;
		Addr <=  "00010010000110";
		Trees_din <= x"0b02880c";
		wait for Clk_period;
		Addr <=  "00010010000111";
		Trees_din <= x"00090508";
		wait for Clk_period;
		Addr <=  "00010010001000";
		Trees_din <= x"00046404";
		wait for Clk_period;
		Addr <=  "00010010001001";
		Trees_din <= x"ffbb1259";
		wait for Clk_period;
		Addr <=  "00010010001010";
		Trees_din <= x"00261259";
		wait for Clk_period;
		Addr <=  "00010010001011";
		Trees_din <= x"ff9f1259";
		wait for Clk_period;
		Addr <=  "00010010001100";
		Trees_din <= x"19008c04";
		wait for Clk_period;
		Addr <=  "00010010001101";
		Trees_din <= x"00641259";
		wait for Clk_period;
		Addr <=  "00010010001110";
		Trees_din <= x"04ff5704";
		wait for Clk_period;
		Addr <=  "00010010001111";
		Trees_din <= x"ffd01259";
		wait for Clk_period;
		Addr <=  "00010010010000";
		Trees_din <= x"002e1259";
		wait for Clk_period;
		Addr <=  "00010010010001";
		Trees_din <= x"1b003a08";
		wait for Clk_period;
		Addr <=  "00010010010010";
		Trees_din <= x"1004c504";
		wait for Clk_period;
		Addr <=  "00010010010011";
		Trees_din <= x"00761259";
		wait for Clk_period;
		Addr <=  "00010010010100";
		Trees_din <= x"001d1259";
		wait for Clk_period;
		Addr <=  "00010010010101";
		Trees_din <= x"ffee1259";
		wait for Clk_period;
		Addr <=  "00010010010110";
		Trees_din <= x"05fc9304";
		wait for Clk_period;
		Addr <=  "00010010010111";
		Trees_din <= x"ff8f12f5";
		wait for Clk_period;
		Addr <=  "00010010011000";
		Trees_din <= x"05005828";
		wait for Clk_period;
		Addr <=  "00010010011001";
		Trees_din <= x"0c008c0c";
		wait for Clk_period;
		Addr <=  "00010010011010";
		Trees_din <= x"01fd4e04";
		wait for Clk_period;
		Addr <=  "00010010011011";
		Trees_din <= x"ffb912f5";
		wait for Clk_period;
		Addr <=  "00010010011100";
		Trees_din <= x"14003304";
		wait for Clk_period;
		Addr <=  "00010010011101";
		Trees_din <= x"ffd812f5";
		wait for Clk_period;
		Addr <=  "00010010011110";
		Trees_din <= x"006912f5";
		wait for Clk_period;
		Addr <=  "00010010011111";
		Trees_din <= x"0700520c";
		wait for Clk_period;
		Addr <=  "00010010100000";
		Trees_din <= x"0b042208";
		wait for Clk_period;
		Addr <=  "00010010100001";
		Trees_din <= x"1a00f304";
		wait for Clk_period;
		Addr <=  "00010010100010";
		Trees_din <= x"007012f5";
		wait for Clk_period;
		Addr <=  "00010010100011";
		Trees_din <= x"ffd612f5";
		wait for Clk_period;
		Addr <=  "00010010100100";
		Trees_din <= x"ffa212f5";
		wait for Clk_period;
		Addr <=  "00010010100101";
		Trees_din <= x"11fd5b08";
		wait for Clk_period;
		Addr <=  "00010010100110";
		Trees_din <= x"19008b04";
		wait for Clk_period;
		Addr <=  "00010010100111";
		Trees_din <= x"004e12f5";
		wait for Clk_period;
		Addr <=  "00010010101000";
		Trees_din <= x"fffe12f5";
		wait for Clk_period;
		Addr <=  "00010010101001";
		Trees_din <= x"06f7f304";
		wait for Clk_period;
		Addr <=  "00010010101010";
		Trees_din <= x"ff7712f5";
		wait for Clk_period;
		Addr <=  "00010010101011";
		Trees_din <= x"ffee12f5";
		wait for Clk_period;
		Addr <=  "00010010101100";
		Trees_din <= x"1202871c";
		wait for Clk_period;
		Addr <=  "00010010101101";
		Trees_din <= x"10046d10";
		wait for Clk_period;
		Addr <=  "00010010101110";
		Trees_din <= x"07005908";
		wait for Clk_period;
		Addr <=  "00010010101111";
		Trees_din <= x"16017e04";
		wait for Clk_period;
		Addr <=  "00010010110000";
		Trees_din <= x"001312f5";
		wait for Clk_period;
		Addr <=  "00010010110001";
		Trees_din <= x"006512f5";
		wait for Clk_period;
		Addr <=  "00010010110010";
		Trees_din <= x"0afedd04";
		wait for Clk_period;
		Addr <=  "00010010110011";
		Trees_din <= x"003d12f5";
		wait for Clk_period;
		Addr <=  "00010010110100";
		Trees_din <= x"ffcf12f5";
		wait for Clk_period;
		Addr <=  "00010010110101";
		Trees_din <= x"05040a08";
		wait for Clk_period;
		Addr <=  "00010010110110";
		Trees_din <= x"03011204";
		wait for Clk_period;
		Addr <=  "00010010110111";
		Trees_din <= x"ff9f12f5";
		wait for Clk_period;
		Addr <=  "00010010111000";
		Trees_din <= x"000e12f5";
		wait for Clk_period;
		Addr <=  "00010010111001";
		Trees_din <= x"003312f5";
		wait for Clk_period;
		Addr <=  "00010010111010";
		Trees_din <= x"10faf604";
		wait for Clk_period;
		Addr <=  "00010010111011";
		Trees_din <= x"001612f5";
		wait for Clk_period;
		Addr <=  "00010010111100";
		Trees_din <= x"ffbc12f5";
		wait for Clk_period;
		Addr <=  "00010010111101";
		Trees_din <= x"05fc9304";
		wait for Clk_period;
		Addr <=  "00010010111110";
		Trees_din <= x"ff921349";
		wait for Clk_period;
		Addr <=  "00010010111111";
		Trees_din <= x"05040a20";
		wait for Clk_period;
		Addr <=  "00010011000000";
		Trees_din <= x"04fbba08";
		wait for Clk_period;
		Addr <=  "00010011000001";
		Trees_din <= x"1d004704";
		wait for Clk_period;
		Addr <=  "00010011000010";
		Trees_din <= x"ff951349";
		wait for Clk_period;
		Addr <=  "00010011000011";
		Trees_din <= x"00041349";
		wait for Clk_period;
		Addr <=  "00010011000100";
		Trees_din <= x"01faee08";
		wait for Clk_period;
		Addr <=  "00010011000101";
		Trees_din <= x"0e010504";
		wait for Clk_period;
		Addr <=  "00010011000110";
		Trees_din <= x"ffa31349";
		wait for Clk_period;
		Addr <=  "00010011000111";
		Trees_din <= x"ffef1349";
		wait for Clk_period;
		Addr <=  "00010011001000";
		Trees_din <= x"07005708";
		wait for Clk_period;
		Addr <=  "00010011001001";
		Trees_din <= x"1400fa04";
		wait for Clk_period;
		Addr <=  "00010011001010";
		Trees_din <= x"003a1349";
		wait for Clk_period;
		Addr <=  "00010011001011";
		Trees_din <= x"fffc1349";
		wait for Clk_period;
		Addr <=  "00010011001100";
		Trees_din <= x"03fe2504";
		wait for Clk_period;
		Addr <=  "00010011001101";
		Trees_din <= x"ff981349";
		wait for Clk_period;
		Addr <=  "00010011001110";
		Trees_din <= x"000d1349";
		wait for Clk_period;
		Addr <=  "00010011001111";
		Trees_din <= x"10027704";
		wait for Clk_period;
		Addr <=  "00010011010000";
		Trees_din <= x"fff91349";
		wait for Clk_period;
		Addr <=  "00010011010001";
		Trees_din <= x"00511349";
		wait for Clk_period;
		Addr <=  "00010011010010";
		Trees_din <= x"05fd6508";
		wait for Clk_period;
		Addr <=  "00010011010011";
		Trees_din <= x"07005004";
		wait for Clk_period;
		Addr <=  "00010011010100";
		Trees_din <= x"002813ad";
		wait for Clk_period;
		Addr <=  "00010011010101";
		Trees_din <= x"ff9313ad";
		wait for Clk_period;
		Addr <=  "00010011010110";
		Trees_din <= x"06f56504";
		wait for Clk_period;
		Addr <=  "00010011010111";
		Trees_din <= x"ffac13ad";
		wait for Clk_period;
		Addr <=  "00010011011000";
		Trees_din <= x"12028718";
		wait for Clk_period;
		Addr <=  "00010011011001";
		Trees_din <= x"01fb1908";
		wait for Clk_period;
		Addr <=  "00010011011010";
		Trees_din <= x"06f9ff04";
		wait for Clk_period;
		Addr <=  "00010011011011";
		Trees_din <= x"ff9f13ad";
		wait for Clk_period;
		Addr <=  "00010011011100";
		Trees_din <= x"001513ad";
		wait for Clk_period;
		Addr <=  "00010011011101";
		Trees_din <= x"0b046808";
		wait for Clk_period;
		Addr <=  "00010011011110";
		Trees_din <= x"0c024e04";
		wait for Clk_period;
		Addr <=  "00010011011111";
		Trees_din <= x"004213ad";
		wait for Clk_period;
		Addr <=  "00010011100000";
		Trees_din <= x"ffef13ad";
		wait for Clk_period;
		Addr <=  "00010011100001";
		Trees_din <= x"19009404";
		wait for Clk_period;
		Addr <=  "00010011100010";
		Trees_din <= x"003e13ad";
		wait for Clk_period;
		Addr <=  "00010011100011";
		Trees_din <= x"ffc113ad";
		wait for Clk_period;
		Addr <=  "00010011100100";
		Trees_din <= x"0f03df0c";
		wait for Clk_period;
		Addr <=  "00010011100101";
		Trees_din <= x"0d03a508";
		wait for Clk_period;
		Addr <=  "00010011100110";
		Trees_din <= x"0501f804";
		wait for Clk_period;
		Addr <=  "00010011100111";
		Trees_din <= x"ff8513ad";
		wait for Clk_period;
		Addr <=  "00010011101000";
		Trees_din <= x"000613ad";
		wait for Clk_period;
		Addr <=  "00010011101001";
		Trees_din <= x"002913ad";
		wait for Clk_period;
		Addr <=  "00010011101010";
		Trees_din <= x"004c13ad";
		wait for Clk_period;
		Addr <=  "00010011101011";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00010011101100";
		Trees_din <= x"05fc9304";
		wait for Clk_period;
		Addr <=  "00010011101101";
		Trees_din <= x"ff9a144d";
		wait for Clk_period;
		Addr <=  "00010011101110";
		Trees_din <= x"0006812c";
		wait for Clk_period;
		Addr <=  "00010011101111";
		Trees_din <= x"0103891c";
		wait for Clk_period;
		Addr <=  "00010011110000";
		Trees_din <= x"05fede0c";
		wait for Clk_period;
		Addr <=  "00010011110001";
		Trees_din <= x"06f76008";
		wait for Clk_period;
		Addr <=  "00010011110010";
		Trees_din <= x"02ffbf04";
		wait for Clk_period;
		Addr <=  "00010011110011";
		Trees_din <= x"0030144d";
		wait for Clk_period;
		Addr <=  "00010011110100";
		Trees_din <= x"ffac144d";
		wait for Clk_period;
		Addr <=  "00010011110101";
		Trees_din <= x"ff97144d";
		wait for Clk_period;
		Addr <=  "00010011110110";
		Trees_din <= x"12007508";
		wait for Clk_period;
		Addr <=  "00010011110111";
		Trees_din <= x"15009e04";
		wait for Clk_period;
		Addr <=  "00010011111000";
		Trees_din <= x"0071144d";
		wait for Clk_period;
		Addr <=  "00010011111001";
		Trees_din <= x"ffe0144d";
		wait for Clk_period;
		Addr <=  "00010011111010";
		Trees_din <= x"0e01bf04";
		wait for Clk_period;
		Addr <=  "00010011111011";
		Trees_din <= x"ffbe144d";
		wait for Clk_period;
		Addr <=  "00010011111100";
		Trees_din <= x"0029144d";
		wait for Clk_period;
		Addr <=  "00010011111101";
		Trees_din <= x"0104bf08";
		wait for Clk_period;
		Addr <=  "00010011111110";
		Trees_din <= x"13ffaf04";
		wait for Clk_period;
		Addr <=  "00010011111111";
		Trees_din <= x"001d144d";
		wait for Clk_period;
		Addr <=  "00010100000000";
		Trees_din <= x"0072144d";
		wait for Clk_period;
		Addr <=  "00010100000001";
		Trees_din <= x"04ffc004";
		wait for Clk_period;
		Addr <=  "00010100000010";
		Trees_din <= x"0040144d";
		wait for Clk_period;
		Addr <=  "00010100000011";
		Trees_din <= x"ffad144d";
		wait for Clk_period;
		Addr <=  "00010100000100";
		Trees_din <= x"0c028618";
		wait for Clk_period;
		Addr <=  "00010100000101";
		Trees_din <= x"07005508";
		wait for Clk_period;
		Addr <=  "00010100000110";
		Trees_din <= x"00090504";
		wait for Clk_period;
		Addr <=  "00010100000111";
		Trees_din <= x"ffee144d";
		wait for Clk_period;
		Addr <=  "00010100001000";
		Trees_din <= x"ffa8144d";
		wait for Clk_period;
		Addr <=  "00010100001001";
		Trees_din <= x"13fdbb08";
		wait for Clk_period;
		Addr <=  "00010100001010";
		Trees_din <= x"05007904";
		wait for Clk_period;
		Addr <=  "00010100001011";
		Trees_din <= x"ffad144d";
		wait for Clk_period;
		Addr <=  "00010100001100";
		Trees_din <= x"001d144d";
		wait for Clk_period;
		Addr <=  "00010100001101";
		Trees_din <= x"1d004204";
		wait for Clk_period;
		Addr <=  "00010100001110";
		Trees_din <= x"fff7144d";
		wait for Clk_period;
		Addr <=  "00010100001111";
		Trees_din <= x"004d144d";
		wait for Clk_period;
		Addr <=  "00010100010000";
		Trees_din <= x"1e005f04";
		wait for Clk_period;
		Addr <=  "00010100010001";
		Trees_din <= x"ffe4144d";
		wait for Clk_period;
		Addr <=  "00010100010010";
		Trees_din <= x"ff99144d";
		wait for Clk_period;
		Addr <=  "00010100010011";
		Trees_din <= x"0500582c";
		wait for Clk_period;
		Addr <=  "00010100010100";
		Trees_din <= x"0004c61c";
		wait for Clk_period;
		Addr <=  "00010100010101";
		Trees_din <= x"0a027614";
		wait for Clk_period;
		Addr <=  "00010100010110";
		Trees_din <= x"1c003a0c";
		wait for Clk_period;
		Addr <=  "00010100010111";
		Trees_din <= x"1e006708";
		wait for Clk_period;
		Addr <=  "00010100011000";
		Trees_din <= x"00025704";
		wait for Clk_period;
		Addr <=  "00010100011001";
		Trees_din <= x"ffd814d9";
		wait for Clk_period;
		Addr <=  "00010100011010";
		Trees_din <= x"003d14d9";
		wait for Clk_period;
		Addr <=  "00010100011011";
		Trees_din <= x"006514d9";
		wait for Clk_period;
		Addr <=  "00010100011100";
		Trees_din <= x"01000404";
		wait for Clk_period;
		Addr <=  "00010100011101";
		Trees_din <= x"ffa614d9";
		wait for Clk_period;
		Addr <=  "00010100011110";
		Trees_din <= x"fff614d9";
		wait for Clk_period;
		Addr <=  "00010100011111";
		Trees_din <= x"01fd6304";
		wait for Clk_period;
		Addr <=  "00010100100000";
		Trees_din <= x"000314d9";
		wait for Clk_period;
		Addr <=  "00010100100001";
		Trees_din <= x"ff9414d9";
		wait for Clk_period;
		Addr <=  "00010100100010";
		Trees_din <= x"0f036108";
		wait for Clk_period;
		Addr <=  "00010100100011";
		Trees_din <= x"0a038904";
		wait for Clk_period;
		Addr <=  "00010100100100";
		Trees_din <= x"ff7f14d9";
		wait for Clk_period;
		Addr <=  "00010100100101";
		Trees_din <= x"001714d9";
		wait for Clk_period;
		Addr <=  "00010100100110";
		Trees_din <= x"13ffcd04";
		wait for Clk_period;
		Addr <=  "00010100100111";
		Trees_din <= x"ffe214d9";
		wait for Clk_period;
		Addr <=  "00010100101000";
		Trees_din <= x"003114d9";
		wait for Clk_period;
		Addr <=  "00010100101001";
		Trees_din <= x"06fa4514";
		wait for Clk_period;
		Addr <=  "00010100101010";
		Trees_din <= x"04ff570c";
		wait for Clk_period;
		Addr <=  "00010100101011";
		Trees_din <= x"19008604";
		wait for Clk_period;
		Addr <=  "00010100101100";
		Trees_din <= x"003414d9";
		wait for Clk_period;
		Addr <=  "00010100101101";
		Trees_din <= x"0e003404";
		wait for Clk_period;
		Addr <=  "00010100101110";
		Trees_din <= x"000414d9";
		wait for Clk_period;
		Addr <=  "00010100101111";
		Trees_din <= x"ffa214d9";
		wait for Clk_period;
		Addr <=  "00010100110000";
		Trees_din <= x"1401bc04";
		wait for Clk_period;
		Addr <=  "00010100110001";
		Trees_din <= x"004f14d9";
		wait for Clk_period;
		Addr <=  "00010100110010";
		Trees_din <= x"fff014d9";
		wait for Clk_period;
		Addr <=  "00010100110011";
		Trees_din <= x"1b003a04";
		wait for Clk_period;
		Addr <=  "00010100110100";
		Trees_din <= x"006114d9";
		wait for Clk_period;
		Addr <=  "00010100110101";
		Trees_din <= x"fff314d9";
		wait for Clk_period;
		Addr <=  "00010100110110";
		Trees_din <= x"05fd6508";
		wait for Clk_period;
		Addr <=  "00010100110111";
		Trees_din <= x"0e03b204";
		wait for Clk_period;
		Addr <=  "00010100111000";
		Trees_din <= x"ff9d1555";
		wait for Clk_period;
		Addr <=  "00010100111001";
		Trees_din <= x"00191555";
		wait for Clk_period;
		Addr <=  "00010100111010";
		Trees_din <= x"06f6be10";
		wait for Clk_period;
		Addr <=  "00010100111011";
		Trees_din <= x"0f005508";
		wait for Clk_period;
		Addr <=  "00010100111100";
		Trees_din <= x"0d032204";
		wait for Clk_period;
		Addr <=  "00010100111101";
		Trees_din <= x"ffdf1555";
		wait for Clk_period;
		Addr <=  "00010100111110";
		Trees_din <= x"00411555";
		wait for Clk_period;
		Addr <=  "00010100111111";
		Trees_din <= x"06f5af04";
		wait for Clk_period;
		Addr <=  "00010101000000";
		Trees_din <= x"ffe31555";
		wait for Clk_period;
		Addr <=  "00010101000001";
		Trees_din <= x"ff9d1555";
		wait for Clk_period;
		Addr <=  "00010101000010";
		Trees_din <= x"0009f01c";
		wait for Clk_period;
		Addr <=  "00010101000011";
		Trees_din <= x"0f015410";
		wait for Clk_period;
		Addr <=  "00010101000100";
		Trees_din <= x"1603d908";
		wait for Clk_period;
		Addr <=  "00010101000101";
		Trees_din <= x"04041b04";
		wait for Clk_period;
		Addr <=  "00010101000110";
		Trees_din <= x"ffb21555";
		wait for Clk_period;
		Addr <=  "00010101000111";
		Trees_din <= x"002b1555";
		wait for Clk_period;
		Addr <=  "00010101001000";
		Trees_din <= x"0f000c04";
		wait for Clk_period;
		Addr <=  "00010101001001";
		Trees_din <= x"ffe71555";
		wait for Clk_period;
		Addr <=  "00010101001010";
		Trees_din <= x"00431555";
		wait for Clk_period;
		Addr <=  "00010101001011";
		Trees_din <= x"18004404";
		wait for Clk_period;
		Addr <=  "00010101001100";
		Trees_din <= x"00631555";
		wait for Clk_period;
		Addr <=  "00010101001101";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00010101001110";
		Trees_din <= x"ffd31555";
		wait for Clk_period;
		Addr <=  "00010101001111";
		Trees_din <= x"001e1555";
		wait for Clk_period;
		Addr <=  "00010101010000";
		Trees_din <= x"0efd8904";
		wait for Clk_period;
		Addr <=  "00010101010001";
		Trees_din <= x"00301555";
		wait for Clk_period;
		Addr <=  "00010101010010";
		Trees_din <= x"04fad304";
		wait for Clk_period;
		Addr <=  "00010101010011";
		Trees_din <= x"fffc1555";
		wait for Clk_period;
		Addr <=  "00010101010100";
		Trees_din <= x"ff981555";
		wait for Clk_period;
		Addr <=  "00010101010101";
		Trees_din <= x"05fec11c";
		wait for Clk_period;
		Addr <=  "00010101010110";
		Trees_din <= x"0e03db14";
		wait for Clk_period;
		Addr <=  "00010101010111";
		Trees_din <= x"00fe2908";
		wait for Clk_period;
		Addr <=  "00010101011000";
		Trees_din <= x"00fce804";
		wait for Clk_period;
		Addr <=  "00010101011001";
		Trees_din <= x"ffcd15d9";
		wait for Clk_period;
		Addr <=  "00010101011010";
		Trees_din <= x"004415d9";
		wait for Clk_period;
		Addr <=  "00010101011011";
		Trees_din <= x"0afabc04";
		wait for Clk_period;
		Addr <=  "00010101011100";
		Trees_din <= x"000715d9";
		wait for Clk_period;
		Addr <=  "00010101011101";
		Trees_din <= x"05fe7004";
		wait for Clk_period;
		Addr <=  "00010101011110";
		Trees_din <= x"ff8015d9";
		wait for Clk_period;
		Addr <=  "00010101011111";
		Trees_din <= x"ffee15d9";
		wait for Clk_period;
		Addr <=  "00010101100000";
		Trees_din <= x"07004f04";
		wait for Clk_period;
		Addr <=  "00010101100001";
		Trees_din <= x"005415d9";
		wait for Clk_period;
		Addr <=  "00010101100010";
		Trees_din <= x"000215d9";
		wait for Clk_period;
		Addr <=  "00010101100011";
		Trees_din <= x"0900510c";
		wait for Clk_period;
		Addr <=  "00010101100100";
		Trees_din <= x"02ffe804";
		wait for Clk_period;
		Addr <=  "00010101100101";
		Trees_din <= x"002715d9";
		wait for Clk_period;
		Addr <=  "00010101100110";
		Trees_din <= x"07005304";
		wait for Clk_period;
		Addr <=  "00010101100111";
		Trees_din <= x"000b15d9";
		wait for Clk_period;
		Addr <=  "00010101101000";
		Trees_din <= x"ffa215d9";
		wait for Clk_period;
		Addr <=  "00010101101001";
		Trees_din <= x"09005408";
		wait for Clk_period;
		Addr <=  "00010101101010";
		Trees_din <= x"0b028704";
		wait for Clk_period;
		Addr <=  "00010101101011";
		Trees_din <= x"005d15d9";
		wait for Clk_period;
		Addr <=  "00010101101100";
		Trees_din <= x"000b15d9";
		wait for Clk_period;
		Addr <=  "00010101101101";
		Trees_din <= x"1d004308";
		wait for Clk_period;
		Addr <=  "00010101101110";
		Trees_din <= x"13001b04";
		wait for Clk_period;
		Addr <=  "00010101101111";
		Trees_din <= x"ffb215d9";
		wait for Clk_period;
		Addr <=  "00010101110000";
		Trees_din <= x"002815d9";
		wait for Clk_period;
		Addr <=  "00010101110001";
		Trees_din <= x"0bfbd604";
		wait for Clk_period;
		Addr <=  "00010101110010";
		Trees_din <= x"ffdb15d9";
		wait for Clk_period;
		Addr <=  "00010101110011";
		Trees_din <= x"0002a804";
		wait for Clk_period;
		Addr <=  "00010101110100";
		Trees_din <= x"005715d9";
		wait for Clk_period;
		Addr <=  "00010101110101";
		Trees_din <= x"000e15d9";
		wait for Clk_period;
		Addr <=  "00010101110110";
		Trees_din <= x"06f50204";
		wait for Clk_period;
		Addr <=  "00010101110111";
		Trees_din <= x"ffa61665";
		wait for Clk_period;
		Addr <=  "00010101111000";
		Trees_din <= x"0500582c";
		wait for Clk_period;
		Addr <=  "00010101111001";
		Trees_din <= x"0c012a14";
		wait for Clk_period;
		Addr <=  "00010101111010";
		Trees_din <= x"0d00bc08";
		wait for Clk_period;
		Addr <=  "00010101111011";
		Trees_din <= x"05ff2604";
		wait for Clk_period;
		Addr <=  "00010101111100";
		Trees_din <= x"ffbd1665";
		wait for Clk_period;
		Addr <=  "00010101111101";
		Trees_din <= x"001e1665";
		wait for Clk_period;
		Addr <=  "00010101111110";
		Trees_din <= x"08006f04";
		wait for Clk_period;
		Addr <=  "00010101111111";
		Trees_din <= x"fff41665";
		wait for Clk_period;
		Addr <=  "00010110000000";
		Trees_din <= x"1700fc04";
		wait for Clk_period;
		Addr <=  "00010110000001";
		Trees_din <= x"00661665";
		wait for Clk_period;
		Addr <=  "00010110000010";
		Trees_din <= x"00101665";
		wait for Clk_period;
		Addr <=  "00010110000011";
		Trees_din <= x"02fe780c";
		wait for Clk_period;
		Addr <=  "00010110000100";
		Trees_din <= x"0a027108";
		wait for Clk_period;
		Addr <=  "00010110000101";
		Trees_din <= x"1d004404";
		wait for Clk_period;
		Addr <=  "00010110000110";
		Trees_din <= x"000e1665";
		wait for Clk_period;
		Addr <=  "00010110000111";
		Trees_din <= x"00501665";
		wait for Clk_period;
		Addr <=  "00010110001000";
		Trees_din <= x"ffad1665";
		wait for Clk_period;
		Addr <=  "00010110001001";
		Trees_din <= x"11fe6004";
		wait for Clk_period;
		Addr <=  "00010110001010";
		Trees_din <= x"00071665";
		wait for Clk_period;
		Addr <=  "00010110001011";
		Trees_din <= x"0d013104";
		wait for Clk_period;
		Addr <=  "00010110001100";
		Trees_din <= x"fff91665";
		wait for Clk_period;
		Addr <=  "00010110001101";
		Trees_din <= x"ff861665";
		wait for Clk_period;
		Addr <=  "00010110001110";
		Trees_din <= x"1300d314";
		wait for Clk_period;
		Addr <=  "00010110001111";
		Trees_din <= x"1004ce0c";
		wait for Clk_period;
		Addr <=  "00010110010000";
		Trees_din <= x"0f036808";
		wait for Clk_period;
		Addr <=  "00010110010001";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00010110010010";
		Trees_din <= x"00111665";
		wait for Clk_period;
		Addr <=  "00010110010011";
		Trees_din <= x"00591665";
		wait for Clk_period;
		Addr <=  "00010110010100";
		Trees_din <= x"ffeb1665";
		wait for Clk_period;
		Addr <=  "00010110010101";
		Trees_din <= x"0f012e04";
		wait for Clk_period;
		Addr <=  "00010110010110";
		Trees_din <= x"ffc81665";
		wait for Clk_period;
		Addr <=  "00010110010111";
		Trees_din <= x"002b1665";
		wait for Clk_period;
		Addr <=  "00010110011000";
		Trees_din <= x"ffdc1665";
		wait for Clk_period;
		Addr <=  "00010110011001";
		Trees_din <= x"05fc9304";
		wait for Clk_period;
		Addr <=  "00010110011010";
		Trees_din <= x"ffaa16b9";
		wait for Clk_period;
		Addr <=  "00010110011011";
		Trees_din <= x"000f0720";
		wait for Clk_period;
		Addr <=  "00010110011100";
		Trees_din <= x"0800660c";
		wait for Clk_period;
		Addr <=  "00010110011101";
		Trees_din <= x"08001708";
		wait for Clk_period;
		Addr <=  "00010110011110";
		Trees_din <= x"17023704";
		wait for Clk_period;
		Addr <=  "00010110011111";
		Trees_din <= x"ffd216b9";
		wait for Clk_period;
		Addr <=  "00010110100000";
		Trees_din <= x"003916b9";
		wait for Clk_period;
		Addr <=  "00010110100001";
		Trees_din <= x"ffb116b9";
		wait for Clk_period;
		Addr <=  "00010110100010";
		Trees_din <= x"1900a70c";
		wait for Clk_period;
		Addr <=  "00010110100011";
		Trees_din <= x"1a00ec08";
		wait for Clk_period;
		Addr <=  "00010110100100";
		Trees_din <= x"1a00a104";
		wait for Clk_period;
		Addr <=  "00010110100101";
		Trees_din <= x"ffdd16b9";
		wait for Clk_period;
		Addr <=  "00010110100110";
		Trees_din <= x"002f16b9";
		wait for Clk_period;
		Addr <=  "00010110100111";
		Trees_din <= x"ffda16b9";
		wait for Clk_period;
		Addr <=  "00010110101000";
		Trees_din <= x"03ff5404";
		wait for Clk_period;
		Addr <=  "00010110101001";
		Trees_din <= x"000816b9";
		wait for Clk_period;
		Addr <=  "00010110101010";
		Trees_din <= x"ffa516b9";
		wait for Clk_period;
		Addr <=  "00010110101011";
		Trees_din <= x"16037404";
		wait for Clk_period;
		Addr <=  "00010110101100";
		Trees_din <= x"ffa816b9";
		wait for Clk_period;
		Addr <=  "00010110101101";
		Trees_din <= x"000a16b9";
		wait for Clk_period;
		Addr <=  "00010110101110";
		Trees_din <= x"05007934";
		wait for Clk_period;
		Addr <=  "00010110101111";
		Trees_din <= x"0c008c10";
		wait for Clk_period;
		Addr <=  "00010110110000";
		Trees_din <= x"0d00bc08";
		wait for Clk_period;
		Addr <=  "00010110110001";
		Trees_din <= x"1c003004";
		wait for Clk_period;
		Addr <=  "00010110110010";
		Trees_din <= x"001a1755";
		wait for Clk_period;
		Addr <=  "00010110110011";
		Trees_din <= x"ffc21755";
		wait for Clk_period;
		Addr <=  "00010110110100";
		Trees_din <= x"10fb2504";
		wait for Clk_period;
		Addr <=  "00010110110101";
		Trees_din <= x"00511755";
		wait for Clk_period;
		Addr <=  "00010110110110";
		Trees_din <= x"00171755";
		wait for Clk_period;
		Addr <=  "00010110110111";
		Trees_din <= x"03041714";
		wait for Clk_period;
		Addr <=  "00010110111000";
		Trees_din <= x"1900920c";
		wait for Clk_period;
		Addr <=  "00010110111001";
		Trees_din <= x"08016d08";
		wait for Clk_period;
		Addr <=  "00010110111010";
		Trees_din <= x"02008604";
		wait for Clk_period;
		Addr <=  "00010110111011";
		Trees_din <= x"ffff1755";
		wait for Clk_period;
		Addr <=  "00010110111100";
		Trees_din <= x"ffad1755";
		wait for Clk_period;
		Addr <=  "00010110111101";
		Trees_din <= x"00391755";
		wait for Clk_period;
		Addr <=  "00010110111110";
		Trees_din <= x"07005104";
		wait for Clk_period;
		Addr <=  "00010110111111";
		Trees_din <= x"ffe21755";
		wait for Clk_period;
		Addr <=  "00010111000000";
		Trees_din <= x"ff851755";
		wait for Clk_period;
		Addr <=  "00010111000001";
		Trees_din <= x"10fb3704";
		wait for Clk_period;
		Addr <=  "00010111000010";
		Trees_din <= x"ffc41755";
		wait for Clk_period;
		Addr <=  "00010111000011";
		Trees_din <= x"01014f08";
		wait for Clk_period;
		Addr <=  "00010111000100";
		Trees_din <= x"14008704";
		wait for Clk_period;
		Addr <=  "00010111000101";
		Trees_din <= x"00301755";
		wait for Clk_period;
		Addr <=  "00010111000110";
		Trees_din <= x"ffd21755";
		wait for Clk_period;
		Addr <=  "00010111000111";
		Trees_din <= x"00551755";
		wait for Clk_period;
		Addr <=  "00010111001000";
		Trees_din <= x"07005810";
		wait for Clk_period;
		Addr <=  "00010111001001";
		Trees_din <= x"14008a04";
		wait for Clk_period;
		Addr <=  "00010111001010";
		Trees_din <= x"ffe51755";
		wait for Clk_period;
		Addr <=  "00010111001011";
		Trees_din <= x"01fb5b04";
		wait for Clk_period;
		Addr <=  "00010111001100";
		Trees_din <= x"fffe1755";
		wait for Clk_period;
		Addr <=  "00010111001101";
		Trees_din <= x"17003204";
		wait for Clk_period;
		Addr <=  "00010111001110";
		Trees_din <= x"00081755";
		wait for Clk_period;
		Addr <=  "00010111001111";
		Trees_din <= x"005e1755";
		wait for Clk_period;
		Addr <=  "00010111010000";
		Trees_din <= x"06fb0208";
		wait for Clk_period;
		Addr <=  "00010111010001";
		Trees_din <= x"06f78904";
		wait for Clk_period;
		Addr <=  "00010111010010";
		Trees_din <= x"00001755";
		wait for Clk_period;
		Addr <=  "00010111010011";
		Trees_din <= x"ffaf1755";
		wait for Clk_period;
		Addr <=  "00010111010100";
		Trees_din <= x"00251755";
		wait for Clk_period;
		Addr <=  "00010111010101";
		Trees_din <= x"00093a30";
		wait for Clk_period;
		Addr <=  "00010111010110";
		Trees_din <= x"06f66f0c";
		wait for Clk_period;
		Addr <=  "00010111010111";
		Trees_din <= x"18004808";
		wait for Clk_period;
		Addr <=  "00010111011000";
		Trees_din <= x"0e026d04";
		wait for Clk_period;
		Addr <=  "00010111011001";
		Trees_din <= x"ffa717d1";
		wait for Clk_period;
		Addr <=  "00010111011010";
		Trees_din <= x"fff517d1";
		wait for Clk_period;
		Addr <=  "00010111011011";
		Trees_din <= x"001717d1";
		wait for Clk_period;
		Addr <=  "00010111011100";
		Trees_din <= x"1a00bf0c";
		wait for Clk_period;
		Addr <=  "00010111011101";
		Trees_din <= x"0afedd04";
		wait for Clk_period;
		Addr <=  "00010111011110";
		Trees_din <= x"ffbe17d1";
		wait for Clk_period;
		Addr <=  "00010111011111";
		Trees_din <= x"00037704";
		wait for Clk_period;
		Addr <=  "00010111100000";
		Trees_din <= x"ffe817d1";
		wait for Clk_period;
		Addr <=  "00010111100001";
		Trees_din <= x"003617d1";
		wait for Clk_period;
		Addr <=  "00010111100010";
		Trees_din <= x"0bfac508";
		wait for Clk_period;
		Addr <=  "00010111100011";
		Trees_din <= x"09005204";
		wait for Clk_period;
		Addr <=  "00010111100100";
		Trees_din <= x"000a17d1";
		wait for Clk_period;
		Addr <=  "00010111100101";
		Trees_din <= x"006e17d1";
		wait for Clk_period;
		Addr <=  "00010111100110";
		Trees_din <= x"1b003608";
		wait for Clk_period;
		Addr <=  "00010111100111";
		Trees_din <= x"0f016804";
		wait for Clk_period;
		Addr <=  "00010111101000";
		Trees_din <= x"ffbb17d1";
		wait for Clk_period;
		Addr <=  "00010111101001";
		Trees_din <= x"001317d1";
		wait for Clk_period;
		Addr <=  "00010111101010";
		Trees_din <= x"1b003904";
		wait for Clk_period;
		Addr <=  "00010111101011";
		Trees_din <= x"005b17d1";
		wait for Clk_period;
		Addr <=  "00010111101100";
		Trees_din <= x"ffe417d1";
		wait for Clk_period;
		Addr <=  "00010111101101";
		Trees_din <= x"0a03890c";
		wait for Clk_period;
		Addr <=  "00010111101110";
		Trees_din <= x"06f94508";
		wait for Clk_period;
		Addr <=  "00010111101111";
		Trees_din <= x"0e003904";
		wait for Clk_period;
		Addr <=  "00010111110000";
		Trees_din <= x"ffe517d1";
		wait for Clk_period;
		Addr <=  "00010111110001";
		Trees_din <= x"ff9e17d1";
		wait for Clk_period;
		Addr <=  "00010111110010";
		Trees_din <= x"fff217d1";
		wait for Clk_period;
		Addr <=  "00010111110011";
		Trees_din <= x"001617d1";
		wait for Clk_period;
		Addr <=  "00010111110100";
		Trees_din <= x"00068128";
		wait for Clk_period;
		Addr <=  "00010111110101";
		Trees_din <= x"01fed914";
		wait for Clk_period;
		Addr <=  "00010111110110";
		Trees_din <= x"0501a40c";
		wait for Clk_period;
		Addr <=  "00010111110111";
		Trees_din <= x"14007204";
		wait for Clk_period;
		Addr <=  "00010111111000";
		Trees_din <= x"0018184d";
		wait for Clk_period;
		Addr <=  "00010111111001";
		Trees_din <= x"10fbfc04";
		wait for Clk_period;
		Addr <=  "00010111111010";
		Trees_din <= x"0009184d";
		wait for Clk_period;
		Addr <=  "00010111111011";
		Trees_din <= x"ff92184d";
		wait for Clk_period;
		Addr <=  "00010111111100";
		Trees_din <= x"02068504";
		wait for Clk_period;
		Addr <=  "00010111111101";
		Trees_din <= x"004a184d";
		wait for Clk_period;
		Addr <=  "00010111111110";
		Trees_din <= x"fff5184d";
		wait for Clk_period;
		Addr <=  "00010111111111";
		Trees_din <= x"05feea0c";
		wait for Clk_period;
		Addr <=  "00011000000000";
		Trees_din <= x"0afabc04";
		wait for Clk_period;
		Addr <=  "00011000000001";
		Trees_din <= x"0034184d";
		wait for Clk_period;
		Addr <=  "00011000000010";
		Trees_din <= x"0f018904";
		wait for Clk_period;
		Addr <=  "00011000000011";
		Trees_din <= x"ffad184d";
		wait for Clk_period;
		Addr <=  "00011000000100";
		Trees_din <= x"0009184d";
		wait for Clk_period;
		Addr <=  "00011000000101";
		Trees_din <= x"06f66904";
		wait for Clk_period;
		Addr <=  "00011000000110";
		Trees_din <= x"0005184d";
		wait for Clk_period;
		Addr <=  "00011000000111";
		Trees_din <= x"004d184d";
		wait for Clk_period;
		Addr <=  "00011000001000";
		Trees_din <= x"0500790c";
		wait for Clk_period;
		Addr <=  "00011000001001";
		Trees_din <= x"1c003604";
		wait for Clk_period;
		Addr <=  "00011000001010";
		Trees_din <= x"ff99184d";
		wait for Clk_period;
		Addr <=  "00011000001011";
		Trees_din <= x"13ffcd04";
		wait for Clk_period;
		Addr <=  "00011000001100";
		Trees_din <= x"ffcf184d";
		wait for Clk_period;
		Addr <=  "00011000001101";
		Trees_din <= x"0020184d";
		wait for Clk_period;
		Addr <=  "00011000001110";
		Trees_din <= x"02060208";
		wait for Clk_period;
		Addr <=  "00011000001111";
		Trees_din <= x"1b003604";
		wait for Clk_period;
		Addr <=  "00011000010000";
		Trees_din <= x"0040184d";
		wait for Clk_period;
		Addr <=  "00011000010001";
		Trees_din <= x"ffed184d";
		wait for Clk_period;
		Addr <=  "00011000010010";
		Trees_din <= x"ffd5184d";
		wait for Clk_period;
		Addr <=  "00011000010011";
		Trees_din <= x"05fd3404";
		wait for Clk_period;
		Addr <=  "00011000010100";
		Trees_din <= x"ffc01899";
		wait for Clk_period;
		Addr <=  "00011000010101";
		Trees_din <= x"11043c20";
		wait for Clk_period;
		Addr <=  "00011000010110";
		Trees_din <= x"0e025f14";
		wait for Clk_period;
		Addr <=  "00011000010111";
		Trees_din <= x"0d037b10";
		wait for Clk_period;
		Addr <=  "00011000011000";
		Trees_din <= x"1b004308";
		wait for Clk_period;
		Addr <=  "00011000011001";
		Trees_din <= x"05040a04";
		wait for Clk_period;
		Addr <=  "00011000011010";
		Trees_din <= x"ffe41899";
		wait for Clk_period;
		Addr <=  "00011000011011";
		Trees_din <= x"00461899";
		wait for Clk_period;
		Addr <=  "00011000011100";
		Trees_din <= x"0b028804";
		wait for Clk_period;
		Addr <=  "00011000011101";
		Trees_din <= x"ffed1899";
		wait for Clk_period;
		Addr <=  "00011000011110";
		Trees_din <= x"00481899";
		wait for Clk_period;
		Addr <=  "00011000011111";
		Trees_din <= x"ffbb1899";
		wait for Clk_period;
		Addr <=  "00011000100000";
		Trees_din <= x"15009e08";
		wait for Clk_period;
		Addr <=  "00011000100001";
		Trees_din <= x"18004304";
		wait for Clk_period;
		Addr <=  "00011000100010";
		Trees_din <= x"00531899";
		wait for Clk_period;
		Addr <=  "00011000100011";
		Trees_din <= x"000c1899";
		wait for Clk_period;
		Addr <=  "00011000100100";
		Trees_din <= x"fff41899";
		wait for Clk_period;
		Addr <=  "00011000100101";
		Trees_din <= x"ffca1899";
		wait for Clk_period;
		Addr <=  "00011000100110";
		Trees_din <= x"0008782c";
		wait for Clk_period;
		Addr <=  "00011000100111";
		Trees_din <= x"05fede10";
		wait for Clk_period;
		Addr <=  "00011000101000";
		Trees_din <= x"0e03db0c";
		wait for Clk_period;
		Addr <=  "00011000101001";
		Trees_din <= x"1900a208";
		wait for Clk_period;
		Addr <=  "00011000101010";
		Trees_din <= x"1b004504";
		wait for Clk_period;
		Addr <=  "00011000101011";
		Trees_din <= x"ff9b1905";
		wait for Clk_period;
		Addr <=  "00011000101100";
		Trees_din <= x"00011905";
		wait for Clk_period;
		Addr <=  "00011000101101";
		Trees_din <= x"00161905";
		wait for Clk_period;
		Addr <=  "00011000101110";
		Trees_din <= x"00351905";
		wait for Clk_period;
		Addr <=  "00011000101111";
		Trees_din <= x"02097618";
		wait for Clk_period;
		Addr <=  "00011000110000";
		Trees_din <= x"03ff7d08";
		wait for Clk_period;
		Addr <=  "00011000110001";
		Trees_din <= x"1003f504";
		wait for Clk_period;
		Addr <=  "00011000110010";
		Trees_din <= x"005b1905";
		wait for Clk_period;
		Addr <=  "00011000110011";
		Trees_din <= x"00011905";
		wait for Clk_period;
		Addr <=  "00011000110100";
		Trees_din <= x"0c010708";
		wait for Clk_period;
		Addr <=  "00011000110101";
		Trees_din <= x"11025d04";
		wait for Clk_period;
		Addr <=  "00011000110110";
		Trees_din <= x"00461905";
		wait for Clk_period;
		Addr <=  "00011000110111";
		Trees_din <= x"00111905";
		wait for Clk_period;
		Addr <=  "00011000111000";
		Trees_din <= x"01ff1e04";
		wait for Clk_period;
		Addr <=  "00011000111001";
		Trees_din <= x"ffc11905";
		wait for Clk_period;
		Addr <=  "00011000111010";
		Trees_din <= x"00151905";
		wait for Clk_period;
		Addr <=  "00011000111011";
		Trees_din <= x"ffd21905";
		wait for Clk_period;
		Addr <=  "00011000111100";
		Trees_din <= x"0a038908";
		wait for Clk_period;
		Addr <=  "00011000111101";
		Trees_din <= x"19008c04";
		wait for Clk_period;
		Addr <=  "00011000111110";
		Trees_din <= x"fffe1905";
		wait for Clk_period;
		Addr <=  "00011000111111";
		Trees_din <= x"ffb11905";
		wait for Clk_period;
		Addr <=  "00011001000000";
		Trees_din <= x"00131905";
		wait for Clk_period;
		Addr <=  "00011001000001";
		Trees_din <= x"05007920";
		wait for Clk_period;
		Addr <=  "00011001000010";
		Trees_din <= x"0c008c08";
		wait for Clk_period;
		Addr <=  "00011001000011";
		Trees_din <= x"0d00bc04";
		wait for Clk_period;
		Addr <=  "00011001000100";
		Trees_din <= x"ffeb1969";
		wait for Clk_period;
		Addr <=  "00011001000101";
		Trees_din <= x"003e1969";
		wait for Clk_period;
		Addr <=  "00011001000110";
		Trees_din <= x"11fe6004";
		wait for Clk_period;
		Addr <=  "00011001000111";
		Trees_din <= x"001b1969";
		wait for Clk_period;
		Addr <=  "00011001001000";
		Trees_din <= x"02ff570c";
		wait for Clk_period;
		Addr <=  "00011001001001";
		Trees_din <= x"0b027508";
		wait for Clk_period;
		Addr <=  "00011001001010";
		Trees_din <= x"07005104";
		wait for Clk_period;
		Addr <=  "00011001001011";
		Trees_din <= x"00461969";
		wait for Clk_period;
		Addr <=  "00011001001100";
		Trees_din <= x"fff61969";
		wait for Clk_period;
		Addr <=  "00011001001101";
		Trees_din <= x"ffc71969";
		wait for Clk_period;
		Addr <=  "00011001001110";
		Trees_din <= x"0b04a504";
		wait for Clk_period;
		Addr <=  "00011001001111";
		Trees_din <= x"ff931969";
		wait for Clk_period;
		Addr <=  "00011001010000";
		Trees_din <= x"ffe61969";
		wait for Clk_period;
		Addr <=  "00011001010001";
		Trees_din <= x"1300d310";
		wait for Clk_period;
		Addr <=  "00011001010010";
		Trees_din <= x"07005808";
		wait for Clk_period;
		Addr <=  "00011001010011";
		Trees_din <= x"1d003e04";
		wait for Clk_period;
		Addr <=  "00011001010100";
		Trees_din <= x"00051969";
		wait for Clk_period;
		Addr <=  "00011001010101";
		Trees_din <= x"004e1969";
		wait for Clk_period;
		Addr <=  "00011001010110";
		Trees_din <= x"07005b04";
		wait for Clk_period;
		Addr <=  "00011001010111";
		Trees_din <= x"ffd71969";
		wait for Clk_period;
		Addr <=  "00011001011000";
		Trees_din <= x"00261969";
		wait for Clk_period;
		Addr <=  "00011001011001";
		Trees_din <= x"ffdf1969";
		wait for Clk_period;
		Addr <=  "00011001011010";
		Trees_din <= x"00068124";
		wait for Clk_period;
		Addr <=  "00011001011011";
		Trees_din <= x"05fede10";
		wait for Clk_period;
		Addr <=  "00011001011100";
		Trees_din <= x"0e03db0c";
		wait for Clk_period;
		Addr <=  "00011001011101";
		Trees_din <= x"07005704";
		wait for Clk_period;
		Addr <=  "00011001011110";
		Trees_din <= x"ffac19cd";
		wait for Clk_period;
		Addr <=  "00011001011111";
		Trees_din <= x"07005804";
		wait for Clk_period;
		Addr <=  "00011001100000";
		Trees_din <= x"003d19cd";
		wait for Clk_period;
		Addr <=  "00011001100001";
		Trees_din <= x"ffd019cd";
		wait for Clk_period;
		Addr <=  "00011001100010";
		Trees_din <= x"003119cd";
		wait for Clk_period;
		Addr <=  "00011001100011";
		Trees_din <= x"0afae904";
		wait for Clk_period;
		Addr <=  "00011001100100";
		Trees_din <= x"ffdf19cd";
		wait for Clk_period;
		Addr <=  "00011001100101";
		Trees_din <= x"1202870c";
		wait for Clk_period;
		Addr <=  "00011001100110";
		Trees_din <= x"1c002d04";
		wait for Clk_period;
		Addr <=  "00011001100111";
		Trees_din <= x"fff519cd";
		wait for Clk_period;
		Addr <=  "00011001101000";
		Trees_din <= x"09005504";
		wait for Clk_period;
		Addr <=  "00011001101001";
		Trees_din <= x"006519cd";
		wait for Clk_period;
		Addr <=  "00011001101010";
		Trees_din <= x"001b19cd";
		wait for Clk_period;
		Addr <=  "00011001101011";
		Trees_din <= x"ffe419cd";
		wait for Clk_period;
		Addr <=  "00011001101100";
		Trees_din <= x"0502b80c";
		wait for Clk_period;
		Addr <=  "00011001101101";
		Trees_din <= x"0d02f208";
		wait for Clk_period;
		Addr <=  "00011001101110";
		Trees_din <= x"1403c904";
		wait for Clk_period;
		Addr <=  "00011001101111";
		Trees_din <= x"ffa019cd";
		wait for Clk_period;
		Addr <=  "00011001110000";
		Trees_din <= x"000b19cd";
		wait for Clk_period;
		Addr <=  "00011001110001";
		Trees_din <= x"000319cd";
		wait for Clk_period;
		Addr <=  "00011001110010";
		Trees_din <= x"001419cd";
		wait for Clk_period;
		Addr <=  "00011001110011";
		Trees_din <= x"1c002204";
		wait for Clk_period;
		Addr <=  "00011001110100";
		Trees_din <= x"002e1a11";
		wait for Clk_period;
		Addr <=  "00011001110101";
		Trees_din <= x"1c002a04";
		wait for Clk_period;
		Addr <=  "00011001110110";
		Trees_din <= x"ffb71a11";
		wait for Clk_period;
		Addr <=  "00011001110111";
		Trees_din <= x"08006808";
		wait for Clk_period;
		Addr <=  "00011001111000";
		Trees_din <= x"0a020f04";
		wait for Clk_period;
		Addr <=  "00011001111001";
		Trees_din <= x"ffad1a11";
		wait for Clk_period;
		Addr <=  "00011001111010";
		Trees_din <= x"00071a11";
		wait for Clk_period;
		Addr <=  "00011001111011";
		Trees_din <= x"08009304";
		wait for Clk_period;
		Addr <=  "00011001111100";
		Trees_din <= x"004a1a11";
		wait for Clk_period;
		Addr <=  "00011001111101";
		Trees_din <= x"0800f008";
		wait for Clk_period;
		Addr <=  "00011001111110";
		Trees_din <= x"09005504";
		wait for Clk_period;
		Addr <=  "00011001111111";
		Trees_din <= x"00031a11";
		wait for Clk_period;
		Addr <=  "00011010000000";
		Trees_din <= x"ffac1a11";
		wait for Clk_period;
		Addr <=  "00011010000001";
		Trees_din <= x"1d003d04";
		wait for Clk_period;
		Addr <=  "00011010000010";
		Trees_din <= x"ffdb1a11";
		wait for Clk_period;
		Addr <=  "00011010000011";
		Trees_din <= x"00201a11";
		wait for Clk_period;
		Addr <=  "00011010000100";
		Trees_din <= x"05005820";
		wait for Clk_period;
		Addr <=  "00011010000101";
		Trees_din <= x"0c008c08";
		wait for Clk_period;
		Addr <=  "00011010000110";
		Trees_din <= x"0d00bc04";
		wait for Clk_period;
		Addr <=  "00011010000111";
		Trees_din <= x"ffee1a75";
		wait for Clk_period;
		Addr <=  "00011010001000";
		Trees_din <= x"00381a75";
		wait for Clk_period;
		Addr <=  "00011010001001";
		Trees_din <= x"07005108";
		wait for Clk_period;
		Addr <=  "00011010001010";
		Trees_din <= x"0e033604";
		wait for Clk_period;
		Addr <=  "00011010001011";
		Trees_din <= x"ffee1a75";
		wait for Clk_period;
		Addr <=  "00011010001100";
		Trees_din <= x"00361a75";
		wait for Clk_period;
		Addr <=  "00011010001101";
		Trees_din <= x"11fd5b04";
		wait for Clk_period;
		Addr <=  "00011010001110";
		Trees_din <= x"001d1a75";
		wait for Clk_period;
		Addr <=  "00011010001111";
		Trees_din <= x"06f7f304";
		wait for Clk_period;
		Addr <=  "00011010010000";
		Trees_din <= x"ff8e1a75";
		wait for Clk_period;
		Addr <=  "00011010010001";
		Trees_din <= x"10041f04";
		wait for Clk_period;
		Addr <=  "00011010010010";
		Trees_din <= x"ffca1a75";
		wait for Clk_period;
		Addr <=  "00011010010011";
		Trees_din <= x"00161a75";
		wait for Clk_period;
		Addr <=  "00011010010100";
		Trees_din <= x"1300d310";
		wait for Clk_period;
		Addr <=  "00011010010101";
		Trees_din <= x"1004ce0c";
		wait for Clk_period;
		Addr <=  "00011010010110";
		Trees_din <= x"06f9ff08";
		wait for Clk_period;
		Addr <=  "00011010010111";
		Trees_din <= x"01fe7c04";
		wait for Clk_period;
		Addr <=  "00011010011000";
		Trees_din <= x"ffe91a75";
		wait for Clk_period;
		Addr <=  "00011010011001";
		Trees_din <= x"00301a75";
		wait for Clk_period;
		Addr <=  "00011010011010";
		Trees_din <= x"004f1a75";
		wait for Clk_period;
		Addr <=  "00011010011011";
		Trees_din <= x"fff41a75";
		wait for Clk_period;
		Addr <=  "00011010011100";
		Trees_din <= x"ffe11a75";
		wait for Clk_period;
		Addr <=  "00011010011101";
		Trees_din <= x"05007920";
		wait for Clk_period;
		Addr <=  "00011010011110";
		Trees_din <= x"0c012a10";
		wait for Clk_period;
		Addr <=  "00011010011111";
		Trees_din <= x"13fd8c04";
		wait for Clk_period;
		Addr <=  "00011010100000";
		Trees_din <= x"ffd51ad1";
		wait for Clk_period;
		Addr <=  "00011010100001";
		Trees_din <= x"0d00a704";
		wait for Clk_period;
		Addr <=  "00011010100010";
		Trees_din <= x"ffee1ad1";
		wait for Clk_period;
		Addr <=  "00011010100011";
		Trees_din <= x"06f7ba04";
		wait for Clk_period;
		Addr <=  "00011010100100";
		Trees_din <= x"00141ad1";
		wait for Clk_period;
		Addr <=  "00011010100101";
		Trees_din <= x"00431ad1";
		wait for Clk_period;
		Addr <=  "00011010100110";
		Trees_din <= x"02fe7808";
		wait for Clk_period;
		Addr <=  "00011010100111";
		Trees_din <= x"1d004404";
		wait for Clk_period;
		Addr <=  "00011010101000";
		Trees_din <= x"ffdc1ad1";
		wait for Clk_period;
		Addr <=  "00011010101001";
		Trees_din <= x"00331ad1";
		wait for Clk_period;
		Addr <=  "00011010101010";
		Trees_din <= x"0d01a304";
		wait for Clk_period;
		Addr <=  "00011010101011";
		Trees_din <= x"fffa1ad1";
		wait for Clk_period;
		Addr <=  "00011010101100";
		Trees_din <= x"ffa41ad1";
		wait for Clk_period;
		Addr <=  "00011010101101";
		Trees_din <= x"0700590c";
		wait for Clk_period;
		Addr <=  "00011010101110";
		Trees_din <= x"0afb1504";
		wait for Clk_period;
		Addr <=  "00011010101111";
		Trees_din <= x"fff11ad1";
		wait for Clk_period;
		Addr <=  "00011010110000";
		Trees_din <= x"09005104";
		wait for Clk_period;
		Addr <=  "00011010110001";
		Trees_din <= x"fffe1ad1";
		wait for Clk_period;
		Addr <=  "00011010110010";
		Trees_din <= x"00491ad1";
		wait for Clk_period;
		Addr <=  "00011010110011";
		Trees_din <= x"ffee1ad1";
		wait for Clk_period;
		Addr <=  "00011010110100";
		Trees_din <= x"00068120";
		wait for Clk_period;
		Addr <=  "00011010110101";
		Trees_din <= x"01fb1904";
		wait for Clk_period;
		Addr <=  "00011010110110";
		Trees_din <= x"ffdd1b2d";
		wait for Clk_period;
		Addr <=  "00011010110111";
		Trees_din <= x"0f001f08";
		wait for Clk_period;
		Addr <=  "00011010111000";
		Trees_din <= x"17027904";
		wait for Clk_period;
		Addr <=  "00011010111001";
		Trees_din <= x"00111b2d";
		wait for Clk_period;
		Addr <=  "00011010111010";
		Trees_din <= x"ffd11b2d";
		wait for Clk_period;
		Addr <=  "00011010111011";
		Trees_din <= x"1102840c";
		wait for Clk_period;
		Addr <=  "00011010111100";
		Trees_din <= x"0d028d08";
		wait for Clk_period;
		Addr <=  "00011010111101";
		Trees_din <= x"1b003704";
		wait for Clk_period;
		Addr <=  "00011010111110";
		Trees_din <= x"00001b2d";
		wait for Clk_period;
		Addr <=  "00011010111111";
		Trees_din <= x"00501b2d";
		wait for Clk_period;
		Addr <=  "00011011000000";
		Trees_din <= x"00021b2d";
		wait for Clk_period;
		Addr <=  "00011011000001";
		Trees_din <= x"1a00d304";
		wait for Clk_period;
		Addr <=  "00011011000010";
		Trees_din <= x"ffd91b2d";
		wait for Clk_period;
		Addr <=  "00011011000011";
		Trees_din <= x"00131b2d";
		wait for Clk_period;
		Addr <=  "00011011000100";
		Trees_din <= x"0c02860c";
		wait for Clk_period;
		Addr <=  "00011011000101";
		Trees_din <= x"07005504";
		wait for Clk_period;
		Addr <=  "00011011000110";
		Trees_din <= x"ffcf1b2d";
		wait for Clk_period;
		Addr <=  "00011011000111";
		Trees_din <= x"07005804";
		wait for Clk_period;
		Addr <=  "00011011001000";
		Trees_din <= x"002d1b2d";
		wait for Clk_period;
		Addr <=  "00011011001001";
		Trees_din <= x"ffeb1b2d";
		wait for Clk_period;
		Addr <=  "00011011001010";
		Trees_din <= x"ffbf1b2d";
		wait for Clk_period;
		Addr <=  "00011011001011";
		Trees_din <= x"0501a424";
		wait for Clk_period;
		Addr <=  "00011011001100";
		Trees_din <= x"1400fa10";
		wait for Clk_period;
		Addr <=  "00011011001101";
		Trees_din <= x"0004c60c";
		wait for Clk_period;
		Addr <=  "00011011001110";
		Trees_din <= x"1a00c304";
		wait for Clk_period;
		Addr <=  "00011011001111";
		Trees_din <= x"fff51b89";
		wait for Clk_period;
		Addr <=  "00011011010000";
		Trees_din <= x"0afca304";
		wait for Clk_period;
		Addr <=  "00011011010001";
		Trees_din <= x"00411b89";
		wait for Clk_period;
		Addr <=  "00011011010010";
		Trees_din <= x"00131b89";
		wait for Clk_period;
		Addr <=  "00011011010011";
		Trees_din <= x"ffdd1b89";
		wait for Clk_period;
		Addr <=  "00011011010100";
		Trees_din <= x"11fd5b04";
		wait for Clk_period;
		Addr <=  "00011011010101";
		Trees_din <= x"001f1b89";
		wait for Clk_period;
		Addr <=  "00011011010110";
		Trees_din <= x"0c008c04";
		wait for Clk_period;
		Addr <=  "00011011010111";
		Trees_din <= x"000f1b89";
		wait for Clk_period;
		Addr <=  "00011011011000";
		Trees_din <= x"0c034208";
		wait for Clk_period;
		Addr <=  "00011011011001";
		Trees_din <= x"19008b04";
		wait for Clk_period;
		Addr <=  "00011011011010";
		Trees_din <= x"ffe41b89";
		wait for Clk_period;
		Addr <=  "00011011011011";
		Trees_din <= x"ff9a1b89";
		wait for Clk_period;
		Addr <=  "00011011011100";
		Trees_din <= x"00031b89";
		wait for Clk_period;
		Addr <=  "00011011011101";
		Trees_din <= x"1601f904";
		wait for Clk_period;
		Addr <=  "00011011011110";
		Trees_din <= x"003d1b89";
		wait for Clk_period;
		Addr <=  "00011011011111";
		Trees_din <= x"0c014c04";
		wait for Clk_period;
		Addr <=  "00011011100000";
		Trees_din <= x"00101b89";
		wait for Clk_period;
		Addr <=  "00011011100001";
		Trees_din <= x"ffdf1b89";
		wait for Clk_period;
		Addr <=  "00011011100010";
		Trees_din <= x"05fec110";
		wait for Clk_period;
		Addr <=  "00011011100011";
		Trees_din <= x"0e03db0c";
		wait for Clk_period;
		Addr <=  "00011011100100";
		Trees_din <= x"00fe2904";
		wait for Clk_period;
		Addr <=  "00011011100101";
		Trees_din <= x"00091bdd";
		wait for Clk_period;
		Addr <=  "00011011100110";
		Trees_din <= x"0bfa2304";
		wait for Clk_period;
		Addr <=  "00011011100111";
		Trees_din <= x"fffa1bdd";
		wait for Clk_period;
		Addr <=  "00011011101000";
		Trees_din <= x"ffa91bdd";
		wait for Clk_period;
		Addr <=  "00011011101001";
		Trees_din <= x"002b1bdd";
		wait for Clk_period;
		Addr <=  "00011011101010";
		Trees_din <= x"04ff5710";
		wait for Clk_period;
		Addr <=  "00011011101011";
		Trees_din <= x"0502b808";
		wait for Clk_period;
		Addr <=  "00011011101100";
		Trees_din <= x"0e003904";
		wait for Clk_period;
		Addr <=  "00011011101101";
		Trees_din <= x"00031bdd";
		wait for Clk_period;
		Addr <=  "00011011101110";
		Trees_din <= x"ffb41bdd";
		wait for Clk_period;
		Addr <=  "00011011101111";
		Trees_din <= x"0800f604";
		wait for Clk_period;
		Addr <=  "00011011110000";
		Trees_din <= x"fff41bdd";
		wait for Clk_period;
		Addr <=  "00011011110001";
		Trees_din <= x"003e1bdd";
		wait for Clk_period;
		Addr <=  "00011011110010";
		Trees_din <= x"0c025b08";
		wait for Clk_period;
		Addr <=  "00011011110011";
		Trees_din <= x"09005104";
		wait for Clk_period;
		Addr <=  "00011011110100";
		Trees_din <= x"fffe1bdd";
		wait for Clk_period;
		Addr <=  "00011011110101";
		Trees_din <= x"003f1bdd";
		wait for Clk_period;
		Addr <=  "00011011110110";
		Trees_din <= x"fff11bdd";
		wait for Clk_period;
		Addr <=  "00011011110111";
		Trees_din <= x"0500791c";
		wait for Clk_period;
		Addr <=  "00011011111000";
		Trees_din <= x"01038910";
		wait for Clk_period;
		Addr <=  "00011011111001";
		Trees_din <= x"11fe6004";
		wait for Clk_period;
		Addr <=  "00011011111010";
		Trees_din <= x"00181c29";
		wait for Clk_period;
		Addr <=  "00011011111011";
		Trees_din <= x"02ff5708";
		wait for Clk_period;
		Addr <=  "00011011111100";
		Trees_din <= x"02fda204";
		wait for Clk_period;
		Addr <=  "00011011111101";
		Trees_din <= x"ffd51c29";
		wait for Clk_period;
		Addr <=  "00011011111110";
		Trees_din <= x"001d1c29";
		wait for Clk_period;
		Addr <=  "00011011111111";
		Trees_din <= x"ffaf1c29";
		wait for Clk_period;
		Addr <=  "00011100000000";
		Trees_din <= x"01063008";
		wait for Clk_period;
		Addr <=  "00011100000001";
		Trees_din <= x"0bfac504";
		wait for Clk_period;
		Addr <=  "00011100000010";
		Trees_din <= x"003c1c29";
		wait for Clk_period;
		Addr <=  "00011100000011";
		Trees_din <= x"000f1c29";
		wait for Clk_period;
		Addr <=  "00011100000100";
		Trees_din <= x"ffe11c29";
		wait for Clk_period;
		Addr <=  "00011100000101";
		Trees_din <= x"07005908";
		wait for Clk_period;
		Addr <=  "00011100000110";
		Trees_din <= x"12020c04";
		wait for Clk_period;
		Addr <=  "00011100000111";
		Trees_din <= x"00371c29";
		wait for Clk_period;
		Addr <=  "00011100001000";
		Trees_din <= x"fffd1c29";
		wait for Clk_period;
		Addr <=  "00011100001001";
		Trees_din <= x"ffef1c29";
		wait for Clk_period;
		Addr <=  "00011100001010";
		Trees_din <= x"05fd3404";
		wait for Clk_period;
		Addr <=  "00011100001011";
		Trees_din <= x"ffd11c6d";
		wait for Clk_period;
		Addr <=  "00011100001100";
		Trees_din <= x"11043c1c";
		wait for Clk_period;
		Addr <=  "00011100001101";
		Trees_din <= x"0e025f14";
		wait for Clk_period;
		Addr <=  "00011100001110";
		Trees_din <= x"05040a10";
		wait for Clk_period;
		Addr <=  "00011100001111";
		Trees_din <= x"0202e708";
		wait for Clk_period;
		Addr <=  "00011100010000";
		Trees_din <= x"09005604";
		wait for Clk_period;
		Addr <=  "00011100010001";
		Trees_din <= x"00221c6d";
		wait for Clk_period;
		Addr <=  "00011100010010";
		Trees_din <= x"ffdc1c6d";
		wait for Clk_period;
		Addr <=  "00011100010011";
		Trees_din <= x"04fee704";
		wait for Clk_period;
		Addr <=  "00011100010100";
		Trees_din <= x"ffbc1c6d";
		wait for Clk_period;
		Addr <=  "00011100010101";
		Trees_din <= x"00071c6d";
		wait for Clk_period;
		Addr <=  "00011100010110";
		Trees_din <= x"002a1c6d";
		wait for Clk_period;
		Addr <=  "00011100010111";
		Trees_din <= x"06f7e504";
		wait for Clk_period;
		Addr <=  "00011100011000";
		Trees_din <= x"00091c6d";
		wait for Clk_period;
		Addr <=  "00011100011001";
		Trees_din <= x"00461c6d";
		wait for Clk_period;
		Addr <=  "00011100011010";
		Trees_din <= x"ffd61c6d";
		wait for Clk_period;
		Addr <=  "00011100011011";
		Trees_din <= x"05fec110";
		wait for Clk_period;
		Addr <=  "00011100011100";
		Trees_din <= x"0e03db0c";
		wait for Clk_period;
		Addr <=  "00011100011101";
		Trees_din <= x"00fe2904";
		wait for Clk_period;
		Addr <=  "00011100011110";
		Trees_din <= x"00081cc1";
		wait for Clk_period;
		Addr <=  "00011100011111";
		Trees_din <= x"0c008904";
		wait for Clk_period;
		Addr <=  "00011100100000";
		Trees_din <= x"fff81cc1";
		wait for Clk_period;
		Addr <=  "00011100100001";
		Trees_din <= x"ffae1cc1";
		wait for Clk_period;
		Addr <=  "00011100100010";
		Trees_din <= x"00281cc1";
		wait for Clk_period;
		Addr <=  "00011100100011";
		Trees_din <= x"09005108";
		wait for Clk_period;
		Addr <=  "00011100100100";
		Trees_din <= x"10044d04";
		wait for Clk_period;
		Addr <=  "00011100100101";
		Trees_din <= x"ffcb1cc1";
		wait for Clk_period;
		Addr <=  "00011100100110";
		Trees_din <= x"000e1cc1";
		wait for Clk_period;
		Addr <=  "00011100100111";
		Trees_din <= x"0009f010";
		wait for Clk_period;
		Addr <=  "00011100101000";
		Trees_din <= x"0c024e0c";
		wait for Clk_period;
		Addr <=  "00011100101001";
		Trees_din <= x"0d02a708";
		wait for Clk_period;
		Addr <=  "00011100101010";
		Trees_din <= x"04014904";
		wait for Clk_period;
		Addr <=  "00011100101011";
		Trees_din <= x"00511cc1";
		wait for Clk_period;
		Addr <=  "00011100101100";
		Trees_din <= x"00171cc1";
		wait for Clk_period;
		Addr <=  "00011100101101";
		Trees_din <= x"00011cc1";
		wait for Clk_period;
		Addr <=  "00011100101110";
		Trees_din <= x"fff91cc1";
		wait for Clk_period;
		Addr <=  "00011100101111";
		Trees_din <= x"ffea1cc1";
		wait for Clk_period;
		Addr <=  "00011100110000";
		Trees_din <= x"04fb5408";
		wait for Clk_period;
		Addr <=  "00011100110001";
		Trees_din <= x"09005504";
		wait for Clk_period;
		Addr <=  "00011100110010";
		Trees_din <= x"ffca1d15";
		wait for Clk_period;
		Addr <=  "00011100110011";
		Trees_din <= x"00061d15";
		wait for Clk_period;
		Addr <=  "00011100110100";
		Trees_din <= x"06f9ff1c";
		wait for Clk_period;
		Addr <=  "00011100110101";
		Trees_din <= x"1e00660c";
		wait for Clk_period;
		Addr <=  "00011100110110";
		Trees_din <= x"01049608";
		wait for Clk_period;
		Addr <=  "00011100110111";
		Trees_din <= x"10fba804";
		wait for Clk_period;
		Addr <=  "00011100111000";
		Trees_din <= x"fffe1d15";
		wait for Clk_period;
		Addr <=  "00011100111001";
		Trees_din <= x"ffb11d15";
		wait for Clk_period;
		Addr <=  "00011100111010";
		Trees_din <= x"00131d15";
		wait for Clk_period;
		Addr <=  "00011100111011";
		Trees_din <= x"1a00c70c";
		wait for Clk_period;
		Addr <=  "00011100111100";
		Trees_din <= x"00feb704";
		wait for Clk_period;
		Addr <=  "00011100111101";
		Trees_din <= x"00221d15";
		wait for Clk_period;
		Addr <=  "00011100111110";
		Trees_din <= x"1d004d04";
		wait for Clk_period;
		Addr <=  "00011100111111";
		Trees_din <= x"ffb51d15";
		wait for Clk_period;
		Addr <=  "00011101000000";
		Trees_din <= x"00011d15";
		wait for Clk_period;
		Addr <=  "00011101000001";
		Trees_din <= x"00421d15";
		wait for Clk_period;
		Addr <=  "00011101000010";
		Trees_din <= x"05001404";
		wait for Clk_period;
		Addr <=  "00011101000011";
		Trees_din <= x"fffd1d15";
		wait for Clk_period;
		Addr <=  "00011101000100";
		Trees_din <= x"00471d15";
		wait for Clk_period;
		Addr <=  "00011101000101";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  6
        -----------
		Addr <=  "00000000000000";
		Trees_din <= x"06091b30";
		wait for Clk_period;
		Addr <=  "00000000000001";
		Trees_din <= x"06054020";
		wait for Clk_period;
		Addr <=  "00000000000010";
		Trees_din <= x"06023214";
		wait for Clk_period;
		Addr <=  "00000000000011";
		Trees_din <= x"06fee904";
		wait for Clk_period;
		Addr <=  "00000000000100";
		Trees_din <= x"ff4d0065";
		wait for Clk_period;
		Addr <=  "00000000000101";
		Trees_din <= x"11fe7f08";
		wait for Clk_period;
		Addr <=  "00000000000110";
		Trees_din <= x"0008bf04";
		wait for Clk_period;
		Addr <=  "00000000000111";
		Trees_din <= x"00b20065";
		wait for Clk_period;
		Addr <=  "00000000001000";
		Trees_din <= x"ff7d0065";
		wait for Clk_period;
		Addr <=  "00000000001001";
		Trees_din <= x"0afae404";
		wait for Clk_period;
		Addr <=  "00000000001010";
		Trees_din <= x"ffe50065";
		wait for Clk_period;
		Addr <=  "00000000001011";
		Trees_din <= x"ff570065";
		wait for Clk_period;
		Addr <=  "00000000001100";
		Trees_din <= x"14010108";
		wait for Clk_period;
		Addr <=  "00000000001101";
		Trees_din <= x"02ffbf04";
		wait for Clk_period;
		Addr <=  "00000000001110";
		Trees_din <= x"013c0065";
		wait for Clk_period;
		Addr <=  "00000000001111";
		Trees_din <= x"ff950065";
		wait for Clk_period;
		Addr <=  "00000000010000";
		Trees_din <= x"ff6b0065";
		wait for Clk_period;
		Addr <=  "00000000010001";
		Trees_din <= x"04f9a008";
		wait for Clk_period;
		Addr <=  "00000000010010";
		Trees_din <= x"09005804";
		wait for Clk_period;
		Addr <=  "00000000010011";
		Trees_din <= x"ff7a0065";
		wait for Clk_period;
		Addr <=  "00000000010100";
		Trees_din <= x"00e20065";
		wait for Clk_period;
		Addr <=  "00000000010101";
		Trees_din <= x"00f95804";
		wait for Clk_period;
		Addr <=  "00000000010110";
		Trees_din <= x"00270065";
		wait for Clk_period;
		Addr <=  "00000000010111";
		Trees_din <= x"02600065";
		wait for Clk_period;
		Addr <=  "00000000011000";
		Trees_din <= x"03d40065";
		wait for Clk_period;
		Addr <=  "00000000011001";
		Trees_din <= x"06054024";
		wait for Clk_period;
		Addr <=  "00000000011010";
		Trees_din <= x"06023218";
		wait for Clk_period;
		Addr <=  "00000000011011";
		Trees_din <= x"06fee904";
		wait for Clk_period;
		Addr <=  "00000000011100";
		Trees_din <= x"ff5400e9";
		wait for Clk_period;
		Addr <=  "00000000011101";
		Trees_din <= x"13f96108";
		wait for Clk_period;
		Addr <=  "00000000011110";
		Trees_din <= x"11fe7f04";
		wait for Clk_period;
		Addr <=  "00000000011111";
		Trees_din <= x"00bc00e9";
		wait for Clk_period;
		Addr <=  "00000000100000";
		Trees_din <= x"ff8700e9";
		wait for Clk_period;
		Addr <=  "00000000100001";
		Trees_din <= x"0afae408";
		wait for Clk_period;
		Addr <=  "00000000100010";
		Trees_din <= x"0003aa04";
		wait for Clk_period;
		Addr <=  "00000000100011";
		Trees_din <= x"003e00e9";
		wait for Clk_period;
		Addr <=  "00000000100100";
		Trees_din <= x"ffa500e9";
		wait for Clk_period;
		Addr <=  "00000000100101";
		Trees_din <= x"ff5d00e9";
		wait for Clk_period;
		Addr <=  "00000000100110";
		Trees_din <= x"0802cf08";
		wait for Clk_period;
		Addr <=  "00000000100111";
		Trees_din <= x"1a00b604";
		wait for Clk_period;
		Addr <=  "00000000101000";
		Trees_din <= x"001e00e9";
		wait for Clk_period;
		Addr <=  "00000000101001";
		Trees_din <= x"ff6f00e9";
		wait for Clk_period;
		Addr <=  "00000000101010";
		Trees_din <= x"00ce00e9";
		wait for Clk_period;
		Addr <=  "00000000101011";
		Trees_din <= x"000a641c";
		wait for Clk_period;
		Addr <=  "00000000101100";
		Trees_din <= x"010c2118";
		wait for Clk_period;
		Addr <=  "00000000101101";
		Trees_din <= x"06091b10";
		wait for Clk_period;
		Addr <=  "00000000101110";
		Trees_din <= x"14014e08";
		wait for Clk_period;
		Addr <=  "00000000101111";
		Trees_din <= x"17006604";
		wait for Clk_period;
		Addr <=  "00000000110000";
		Trees_din <= x"003a00e9";
		wait for Clk_period;
		Addr <=  "00000000110001";
		Trees_din <= x"ff9000e9";
		wait for Clk_period;
		Addr <=  "00000000110010";
		Trees_din <= x"11ff2e04";
		wait for Clk_period;
		Addr <=  "00000000110011";
		Trees_din <= x"ff9f00e9";
		wait for Clk_period;
		Addr <=  "00000000110100";
		Trees_din <= x"01f700e9";
		wait for Clk_period;
		Addr <=  "00000000110101";
		Trees_din <= x"13025704";
		wait for Clk_period;
		Addr <=  "00000000110110";
		Trees_din <= x"01c100e9";
		wait for Clk_period;
		Addr <=  "00000000110111";
		Trees_din <= x"008b00e9";
		wait for Clk_period;
		Addr <=  "00000000111000";
		Trees_din <= x"ffa000e9";
		wait for Clk_period;
		Addr <=  "00000000111001";
		Trees_din <= x"ff8500e9";
		wait for Clk_period;
		Addr <=  "00000000111010";
		Trees_din <= x"0605401c";
		wait for Clk_period;
		Addr <=  "00000000111011";
		Trees_din <= x"06fee904";
		wait for Clk_period;
		Addr <=  "00000000111100";
		Trees_din <= x"ff580155";
		wait for Clk_period;
		Addr <=  "00000000111101";
		Trees_din <= x"13f9610c";
		wait for Clk_period;
		Addr <=  "00000000111110";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00000000111111";
		Trees_din <= x"013d0155";
		wait for Clk_period;
		Addr <=  "00000001000000";
		Trees_din <= x"12fe6204";
		wait for Clk_period;
		Addr <=  "00000001000001";
		Trees_din <= x"00380155";
		wait for Clk_period;
		Addr <=  "00000001000010";
		Trees_din <= x"ff850155";
		wait for Clk_period;
		Addr <=  "00000001000011";
		Trees_din <= x"0afae408";
		wait for Clk_period;
		Addr <=  "00000001000100";
		Trees_din <= x"18004304";
		wait for Clk_period;
		Addr <=  "00000001000101";
		Trees_din <= x"ff870155";
		wait for Clk_period;
		Addr <=  "00000001000110";
		Trees_din <= x"00ce0155";
		wait for Clk_period;
		Addr <=  "00000001000111";
		Trees_din <= x"ff600155";
		wait for Clk_period;
		Addr <=  "00000001001000";
		Trees_din <= x"000a6418";
		wait for Clk_period;
		Addr <=  "00000001001001";
		Trees_din <= x"01070110";
		wait for Clk_period;
		Addr <=  "00000001001010";
		Trees_din <= x"06091b0c";
		wait for Clk_period;
		Addr <=  "00000001001011";
		Trees_din <= x"0308a908";
		wait for Clk_period;
		Addr <=  "00000001001100";
		Trees_din <= x"0b028804";
		wait for Clk_period;
		Addr <=  "00000001001101";
		Trees_din <= x"014c0155";
		wait for Clk_period;
		Addr <=  "00000001001110";
		Trees_din <= x"fff60155";
		wait for Clk_period;
		Addr <=  "00000001001111";
		Trees_din <= x"ff9e0155";
		wait for Clk_period;
		Addr <=  "00000001010000";
		Trees_din <= x"013f0155";
		wait for Clk_period;
		Addr <=  "00000001010001";
		Trees_din <= x"17000004";
		wait for Clk_period;
		Addr <=  "00000001010010";
		Trees_din <= x"00e20155";
		wait for Clk_period;
		Addr <=  "00000001010011";
		Trees_din <= x"ff850155";
		wait for Clk_period;
		Addr <=  "00000001010100";
		Trees_din <= x"ff8e0155";
		wait for Clk_period;
		Addr <=  "00000001010101";
		Trees_din <= x"0605401c";
		wait for Clk_period;
		Addr <=  "00000001010110";
		Trees_din <= x"06fee904";
		wait for Clk_period;
		Addr <=  "00000001010111";
		Trees_din <= x"ff5b01c9";
		wait for Clk_period;
		Addr <=  "00000001011000";
		Trees_din <= x"13f9610c";
		wait for Clk_period;
		Addr <=  "00000001011001";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00000001011010";
		Trees_din <= x"010401c9";
		wait for Clk_period;
		Addr <=  "00000001011011";
		Trees_din <= x"07005704";
		wait for Clk_period;
		Addr <=  "00000001011100";
		Trees_din <= x"003701c9";
		wait for Clk_period;
		Addr <=  "00000001011101";
		Trees_din <= x"ff8c01c9";
		wait for Clk_period;
		Addr <=  "00000001011110";
		Trees_din <= x"0afae408";
		wait for Clk_period;
		Addr <=  "00000001011111";
		Trees_din <= x"18004304";
		wait for Clk_period;
		Addr <=  "00000001100000";
		Trees_din <= x"ff8c01c9";
		wait for Clk_period;
		Addr <=  "00000001100001";
		Trees_din <= x"00ae01c9";
		wait for Clk_period;
		Addr <=  "00000001100010";
		Trees_din <= x"ff6401c9";
		wait for Clk_period;
		Addr <=  "00000001100011";
		Trees_din <= x"000a641c";
		wait for Clk_period;
		Addr <=  "00000001100100";
		Trees_din <= x"02026c10";
		wait for Clk_period;
		Addr <=  "00000001100101";
		Trees_din <= x"13019608";
		wait for Clk_period;
		Addr <=  "00000001100110";
		Trees_din <= x"11fd0404";
		wait for Clk_period;
		Addr <=  "00000001100111";
		Trees_din <= x"005301c9";
		wait for Clk_period;
		Addr <=  "00000001101000";
		Trees_din <= x"010201c9";
		wait for Clk_period;
		Addr <=  "00000001101001";
		Trees_din <= x"06103104";
		wait for Clk_period;
		Addr <=  "00000001101010";
		Trees_din <= x"ff9801c9";
		wait for Clk_period;
		Addr <=  "00000001101011";
		Trees_din <= x"00bc01c9";
		wait for Clk_period;
		Addr <=  "00000001101100";
		Trees_din <= x"19007904";
		wait for Clk_period;
		Addr <=  "00000001101101";
		Trees_din <= x"00a401c9";
		wait for Clk_period;
		Addr <=  "00000001101110";
		Trees_din <= x"17006604";
		wait for Clk_period;
		Addr <=  "00000001101111";
		Trees_din <= x"001101c9";
		wait for Clk_period;
		Addr <=  "00000001110000";
		Trees_din <= x"ff9b01c9";
		wait for Clk_period;
		Addr <=  "00000001110001";
		Trees_din <= x"ff9601c9";
		wait for Clk_period;
		Addr <=  "00000001110010";
		Trees_din <= x"06054024";
		wait for Clk_period;
		Addr <=  "00000001110011";
		Trees_din <= x"06fee90c";
		wait for Clk_period;
		Addr <=  "00000001110100";
		Trees_din <= x"1703fd04";
		wait for Clk_period;
		Addr <=  "00000001110101";
		Trees_din <= x"ff5e024d";
		wait for Clk_period;
		Addr <=  "00000001110110";
		Trees_din <= x"10042704";
		wait for Clk_period;
		Addr <=  "00000001110111";
		Trees_din <= x"ff7a024d";
		wait for Clk_period;
		Addr <=  "00000001111000";
		Trees_din <= x"0038024d";
		wait for Clk_period;
		Addr <=  "00000001111001";
		Trees_din <= x"13f9610c";
		wait for Clk_period;
		Addr <=  "00000001111010";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00000001111011";
		Trees_din <= x"00e2024d";
		wait for Clk_period;
		Addr <=  "00000001111100";
		Trees_din <= x"11fe7f04";
		wait for Clk_period;
		Addr <=  "00000001111101";
		Trees_din <= x"003b024d";
		wait for Clk_period;
		Addr <=  "00000001111110";
		Trees_din <= x"ff91024d";
		wait for Clk_period;
		Addr <=  "00000001111111";
		Trees_din <= x"0afae408";
		wait for Clk_period;
		Addr <=  "00000010000000";
		Trees_din <= x"18004304";
		wait for Clk_period;
		Addr <=  "00000010000001";
		Trees_din <= x"ff92024d";
		wait for Clk_period;
		Addr <=  "00000010000010";
		Trees_din <= x"0098024d";
		wait for Clk_period;
		Addr <=  "00000010000011";
		Trees_din <= x"ff69024d";
		wait for Clk_period;
		Addr <=  "00000010000100";
		Trees_din <= x"000a641c";
		wait for Clk_period;
		Addr <=  "00000010000101";
		Trees_din <= x"06091b14";
		wait for Clk_period;
		Addr <=  "00000010000110";
		Trees_din <= x"0b02880c";
		wait for Clk_period;
		Addr <=  "00000010000111";
		Trees_din <= x"14014e04";
		wait for Clk_period;
		Addr <=  "00000010001000";
		Trees_din <= x"fff0024d";
		wait for Clk_period;
		Addr <=  "00000010001001";
		Trees_din <= x"00f9b904";
		wait for Clk_period;
		Addr <=  "00000010001010";
		Trees_din <= x"0026024d";
		wait for Clk_period;
		Addr <=  "00000010001011";
		Trees_din <= x"00ed024d";
		wait for Clk_period;
		Addr <=  "00000010001100";
		Trees_din <= x"03fb7404";
		wait for Clk_period;
		Addr <=  "00000010001101";
		Trees_din <= x"0021024d";
		wait for Clk_period;
		Addr <=  "00000010001110";
		Trees_din <= x"ff89024d";
		wait for Clk_period;
		Addr <=  "00000010001111";
		Trees_din <= x"13025704";
		wait for Clk_period;
		Addr <=  "00000010010000";
		Trees_din <= x"00e2024d";
		wait for Clk_period;
		Addr <=  "00000010010001";
		Trees_din <= x"004d024d";
		wait for Clk_period;
		Addr <=  "00000010010010";
		Trees_din <= x"ff9f024d";
		wait for Clk_period;
		Addr <=  "00000010010011";
		Trees_din <= x"06054024";
		wait for Clk_period;
		Addr <=  "00000010010100";
		Trees_din <= x"06fee90c";
		wait for Clk_period;
		Addr <=  "00000010010101";
		Trees_din <= x"1703fd04";
		wait for Clk_period;
		Addr <=  "00000010010110";
		Trees_din <= x"ff6002d9";
		wait for Clk_period;
		Addr <=  "00000010010111";
		Trees_din <= x"04012004";
		wait for Clk_period;
		Addr <=  "00000010011000";
		Trees_din <= x"ff8002d9";
		wait for Clk_period;
		Addr <=  "00000010011001";
		Trees_din <= x"003d02d9";
		wait for Clk_period;
		Addr <=  "00000010011010";
		Trees_din <= x"13f9610c";
		wait for Clk_period;
		Addr <=  "00000010011011";
		Trees_din <= x"07005808";
		wait for Clk_period;
		Addr <=  "00000010011100";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00000010011101";
		Trees_din <= x"00e902d9";
		wait for Clk_period;
		Addr <=  "00000010011110";
		Trees_din <= x"001502d9";
		wait for Clk_period;
		Addr <=  "00000010011111";
		Trees_din <= x"ff9902d9";
		wait for Clk_period;
		Addr <=  "00000010100000";
		Trees_din <= x"0afae408";
		wait for Clk_period;
		Addr <=  "00000010100001";
		Trees_din <= x"18004304";
		wait for Clk_period;
		Addr <=  "00000010100010";
		Trees_din <= x"ff9702d9";
		wait for Clk_period;
		Addr <=  "00000010100011";
		Trees_din <= x"008402d9";
		wait for Clk_period;
		Addr <=  "00000010100100";
		Trees_din <= x"ff6d02d9";
		wait for Clk_period;
		Addr <=  "00000010100101";
		Trees_din <= x"06091b14";
		wait for Clk_period;
		Addr <=  "00000010100110";
		Trees_din <= x"14014e08";
		wait for Clk_period;
		Addr <=  "00000010100111";
		Trees_din <= x"1900a004";
		wait for Clk_period;
		Addr <=  "00000010101000";
		Trees_din <= x"ff8702d9";
		wait for Clk_period;
		Addr <=  "00000010101001";
		Trees_din <= x"001702d9";
		wait for Clk_period;
		Addr <=  "00000010101010";
		Trees_din <= x"11ff2e04";
		wait for Clk_period;
		Addr <=  "00000010101011";
		Trees_din <= x"ffa602d9";
		wait for Clk_period;
		Addr <=  "00000010101100";
		Trees_din <= x"07005a04";
		wait for Clk_period;
		Addr <=  "00000010101101";
		Trees_din <= x"00c302d9";
		wait for Clk_period;
		Addr <=  "00000010101110";
		Trees_din <= x"001402d9";
		wait for Clk_period;
		Addr <=  "00000010101111";
		Trees_din <= x"0201540c";
		wait for Clk_period;
		Addr <=  "00000010110000";
		Trees_din <= x"13025708";
		wait for Clk_period;
		Addr <=  "00000010110001";
		Trees_din <= x"15007604";
		wait for Clk_period;
		Addr <=  "00000010110010";
		Trees_din <= x"003902d9";
		wait for Clk_period;
		Addr <=  "00000010110011";
		Trees_din <= x"00cf02d9";
		wait for Clk_period;
		Addr <=  "00000010110100";
		Trees_din <= x"004102d9";
		wait for Clk_period;
		Addr <=  "00000010110101";
		Trees_din <= x"002a02d9";
		wait for Clk_period;
		Addr <=  "00000010110110";
		Trees_din <= x"06054020";
		wait for Clk_period;
		Addr <=  "00000010110111";
		Trees_din <= x"06fee90c";
		wait for Clk_period;
		Addr <=  "00000010111000";
		Trees_din <= x"1703fd04";
		wait for Clk_period;
		Addr <=  "00000010111001";
		Trees_din <= x"ff610365";
		wait for Clk_period;
		Addr <=  "00000010111010";
		Trees_din <= x"0f000804";
		wait for Clk_period;
		Addr <=  "00000010111011";
		Trees_din <= x"ff870365";
		wait for Clk_period;
		Addr <=  "00000010111100";
		Trees_din <= x"00390365";
		wait for Clk_period;
		Addr <=  "00000010111101";
		Trees_din <= x"13ff6710";
		wait for Clk_period;
		Addr <=  "00000010111110";
		Trees_din <= x"0c02cf08";
		wait for Clk_period;
		Addr <=  "00000010111111";
		Trees_din <= x"04fccf04";
		wait for Clk_period;
		Addr <=  "00000011000000";
		Trees_din <= x"ff7e0365";
		wait for Clk_period;
		Addr <=  "00000011000001";
		Trees_din <= x"00770365";
		wait for Clk_period;
		Addr <=  "00000011000010";
		Trees_din <= x"05fbd404";
		wait for Clk_period;
		Addr <=  "00000011000011";
		Trees_din <= x"ffff0365";
		wait for Clk_period;
		Addr <=  "00000011000100";
		Trees_din <= x"00d40365";
		wait for Clk_period;
		Addr <=  "00000011000101";
		Trees_din <= x"ff730365";
		wait for Clk_period;
		Addr <=  "00000011000110";
		Trees_din <= x"06091b18";
		wait for Clk_period;
		Addr <=  "00000011000111";
		Trees_din <= x"0b028810";
		wait for Clk_period;
		Addr <=  "00000011001000";
		Trees_din <= x"07005908";
		wait for Clk_period;
		Addr <=  "00000011001001";
		Trees_din <= x"09005504";
		wait for Clk_period;
		Addr <=  "00000011001010";
		Trees_din <= x"fff60365";
		wait for Clk_period;
		Addr <=  "00000011001011";
		Trees_din <= x"00c80365";
		wait for Clk_period;
		Addr <=  "00000011001100";
		Trees_din <= x"01ffc504";
		wait for Clk_period;
		Addr <=  "00000011001101";
		Trees_din <= x"00140365";
		wait for Clk_period;
		Addr <=  "00000011001110";
		Trees_din <= x"ffe60365";
		wait for Clk_period;
		Addr <=  "00000011001111";
		Trees_din <= x"03fa5a04";
		wait for Clk_period;
		Addr <=  "00000011010000";
		Trees_din <= x"00130365";
		wait for Clk_period;
		Addr <=  "00000011010001";
		Trees_din <= x"ff8e0365";
		wait for Clk_period;
		Addr <=  "00000011010010";
		Trees_din <= x"03f59204";
		wait for Clk_period;
		Addr <=  "00000011010011";
		Trees_din <= x"001a0365";
		wait for Clk_period;
		Addr <=  "00000011010100";
		Trees_din <= x"13025708";
		wait for Clk_period;
		Addr <=  "00000011010101";
		Trees_din <= x"07004e04";
		wait for Clk_period;
		Addr <=  "00000011010110";
		Trees_din <= x"00430365";
		wait for Clk_period;
		Addr <=  "00000011010111";
		Trees_din <= x"00c20365";
		wait for Clk_period;
		Addr <=  "00000011011000";
		Trees_din <= x"00360365";
		wait for Clk_period;
		Addr <=  "00000011011001";
		Trees_din <= x"0602321c";
		wait for Clk_period;
		Addr <=  "00000011011010";
		Trees_din <= x"06fee90c";
		wait for Clk_period;
		Addr <=  "00000011011011";
		Trees_din <= x"1703fd04";
		wait for Clk_period;
		Addr <=  "00000011011100";
		Trees_din <= x"ff6203d9";
		wait for Clk_period;
		Addr <=  "00000011011101";
		Trees_din <= x"0303cb04";
		wait for Clk_period;
		Addr <=  "00000011011110";
		Trees_din <= x"ff8d03d9";
		wait for Clk_period;
		Addr <=  "00000011011111";
		Trees_din <= x"004203d9";
		wait for Clk_period;
		Addr <=  "00000011100000";
		Trees_din <= x"1201910c";
		wait for Clk_period;
		Addr <=  "00000011100001";
		Trees_din <= x"0003aa08";
		wait for Clk_period;
		Addr <=  "00000011100010";
		Trees_din <= x"11fe7f04";
		wait for Clk_period;
		Addr <=  "00000011100011";
		Trees_din <= x"00aa03d9";
		wait for Clk_period;
		Addr <=  "00000011100100";
		Trees_din <= x"002103d9";
		wait for Clk_period;
		Addr <=  "00000011100101";
		Trees_din <= x"ff9503d9";
		wait for Clk_period;
		Addr <=  "00000011100110";
		Trees_din <= x"ff7a03d9";
		wait for Clk_period;
		Addr <=  "00000011100111";
		Trees_din <= x"06091b14";
		wait for Clk_period;
		Addr <=  "00000011101000";
		Trees_din <= x"0b047410";
		wait for Clk_period;
		Addr <=  "00000011101001";
		Trees_din <= x"0105950c";
		wait for Clk_period;
		Addr <=  "00000011101010";
		Trees_din <= x"01fac304";
		wait for Clk_period;
		Addr <=  "00000011101011";
		Trees_din <= x"ffa703d9";
		wait for Clk_period;
		Addr <=  "00000011101100";
		Trees_din <= x"0c009904";
		wait for Clk_period;
		Addr <=  "00000011101101";
		Trees_din <= x"fff903d9";
		wait for Clk_period;
		Addr <=  "00000011101110";
		Trees_din <= x"00b103d9";
		wait for Clk_period;
		Addr <=  "00000011101111";
		Trees_din <= x"ffa403d9";
		wait for Clk_period;
		Addr <=  "00000011110000";
		Trees_din <= x"ff9003d9";
		wait for Clk_period;
		Addr <=  "00000011110001";
		Trees_din <= x"0bfacb08";
		wait for Clk_period;
		Addr <=  "00000011110010";
		Trees_din <= x"06103104";
		wait for Clk_period;
		Addr <=  "00000011110011";
		Trees_din <= x"ffb403d9";
		wait for Clk_period;
		Addr <=  "00000011110100";
		Trees_din <= x"009503d9";
		wait for Clk_period;
		Addr <=  "00000011110101";
		Trees_din <= x"00b803d9";
		wait for Clk_period;
		Addr <=  "00000011110110";
		Trees_din <= x"0602321c";
		wait for Clk_period;
		Addr <=  "00000011110111";
		Trees_din <= x"06fee90c";
		wait for Clk_period;
		Addr <=  "00000011111000";
		Trees_din <= x"1703fd04";
		wait for Clk_period;
		Addr <=  "00000011111001";
		Trees_din <= x"ff630455";
		wait for Clk_period;
		Addr <=  "00000011111010";
		Trees_din <= x"0f000804";
		wait for Clk_period;
		Addr <=  "00000011111011";
		Trees_din <= x"ff930455";
		wait for Clk_period;
		Addr <=  "00000011111100";
		Trees_din <= x"00470455";
		wait for Clk_period;
		Addr <=  "00000011111101";
		Trees_din <= x"1201910c";
		wait for Clk_period;
		Addr <=  "00000011111110";
		Trees_din <= x"0003aa08";
		wait for Clk_period;
		Addr <=  "00000011111111";
		Trees_din <= x"11fe7f04";
		wait for Clk_period;
		Addr <=  "00000100000000";
		Trees_din <= x"00980455";
		wait for Clk_period;
		Addr <=  "00000100000001";
		Trees_din <= x"001f0455";
		wait for Clk_period;
		Addr <=  "00000100000010";
		Trees_din <= x"ff9c0455";
		wait for Clk_period;
		Addr <=  "00000100000011";
		Trees_din <= x"ff7e0455";
		wait for Clk_period;
		Addr <=  "00000100000100";
		Trees_din <= x"06091b18";
		wait for Clk_period;
		Addr <=  "00000100000101";
		Trees_din <= x"0b047414";
		wait for Clk_period;
		Addr <=  "00000100000110";
		Trees_din <= x"04f9a00c";
		wait for Clk_period;
		Addr <=  "00000100000111";
		Trees_din <= x"12020004";
		wait for Clk_period;
		Addr <=  "00000100001000";
		Trees_din <= x"ff7f0455";
		wait for Clk_period;
		Addr <=  "00000100001001";
		Trees_din <= x"17000004";
		wait for Clk_period;
		Addr <=  "00000100001010";
		Trees_din <= x"00970455";
		wait for Clk_period;
		Addr <=  "00000100001011";
		Trees_din <= x"fffc0455";
		wait for Clk_period;
		Addr <=  "00000100001100";
		Trees_din <= x"0bfabb04";
		wait for Clk_period;
		Addr <=  "00000100001101";
		Trees_din <= x"fffc0455";
		wait for Clk_period;
		Addr <=  "00000100001110";
		Trees_din <= x"009b0455";
		wait for Clk_period;
		Addr <=  "00000100001111";
		Trees_din <= x"ff950455";
		wait for Clk_period;
		Addr <=  "00000100010000";
		Trees_din <= x"0bfacb08";
		wait for Clk_period;
		Addr <=  "00000100010001";
		Trees_din <= x"06103104";
		wait for Clk_period;
		Addr <=  "00000100010010";
		Trees_din <= x"ffb90455";
		wait for Clk_period;
		Addr <=  "00000100010011";
		Trees_din <= x"008a0455";
		wait for Clk_period;
		Addr <=  "00000100010100";
		Trees_din <= x"00b00455";
		wait for Clk_period;
		Addr <=  "00000100010101";
		Trees_din <= x"0602321c";
		wait for Clk_period;
		Addr <=  "00000100010110";
		Trees_din <= x"06fee90c";
		wait for Clk_period;
		Addr <=  "00000100010111";
		Trees_din <= x"16040004";
		wait for Clk_period;
		Addr <=  "00000100011000";
		Trees_din <= x"ff6404d1";
		wait for Clk_period;
		Addr <=  "00000100011001";
		Trees_din <= x"19009004";
		wait for Clk_period;
		Addr <=  "00000100011010";
		Trees_din <= x"ff9c04d1";
		wait for Clk_period;
		Addr <=  "00000100011011";
		Trees_din <= x"004804d1";
		wait for Clk_period;
		Addr <=  "00000100011100";
		Trees_din <= x"1201910c";
		wait for Clk_period;
		Addr <=  "00000100011101";
		Trees_din <= x"0003aa08";
		wait for Clk_period;
		Addr <=  "00000100011110";
		Trees_din <= x"03fbbc04";
		wait for Clk_period;
		Addr <=  "00000100011111";
		Trees_din <= x"009204d1";
		wait for Clk_period;
		Addr <=  "00000100100000";
		Trees_din <= x"001204d1";
		wait for Clk_period;
		Addr <=  "00000100100001";
		Trees_din <= x"ffa204d1";
		wait for Clk_period;
		Addr <=  "00000100100010";
		Trees_din <= x"ff8304d1";
		wait for Clk_period;
		Addr <=  "00000100100011";
		Trees_din <= x"06091b18";
		wait for Clk_period;
		Addr <=  "00000100100100";
		Trees_din <= x"0b047414";
		wait for Clk_period;
		Addr <=  "00000100100101";
		Trees_din <= x"01059510";
		wait for Clk_period;
		Addr <=  "00000100100110";
		Trees_din <= x"12020008";
		wait for Clk_period;
		Addr <=  "00000100100111";
		Trees_din <= x"04f9a004";
		wait for Clk_period;
		Addr <=  "00000100101000";
		Trees_din <= x"ff8a04d1";
		wait for Clk_period;
		Addr <=  "00000100101001";
		Trees_din <= x"007304d1";
		wait for Clk_period;
		Addr <=  "00000100101010";
		Trees_din <= x"09005604";
		wait for Clk_period;
		Addr <=  "00000100101011";
		Trees_din <= x"001d04d1";
		wait for Clk_period;
		Addr <=  "00000100101100";
		Trees_din <= x"00a604d1";
		wait for Clk_period;
		Addr <=  "00000100101101";
		Trees_din <= x"ffab04d1";
		wait for Clk_period;
		Addr <=  "00000100101110";
		Trees_din <= x"ff9a04d1";
		wait for Clk_period;
		Addr <=  "00000100101111";
		Trees_din <= x"0bfacb08";
		wait for Clk_period;
		Addr <=  "00000100110000";
		Trees_din <= x"06103104";
		wait for Clk_period;
		Addr <=  "00000100110001";
		Trees_din <= x"ffbd04d1";
		wait for Clk_period;
		Addr <=  "00000100110010";
		Trees_din <= x"008004d1";
		wait for Clk_period;
		Addr <=  "00000100110011";
		Trees_din <= x"00a904d1";
		wait for Clk_period;
		Addr <=  "00000100110100";
		Trees_din <= x"0602321c";
		wait for Clk_period;
		Addr <=  "00000100110101";
		Trees_din <= x"06fee90c";
		wait for Clk_period;
		Addr <=  "00000100110110";
		Trees_din <= x"1703fd04";
		wait for Clk_period;
		Addr <=  "00000100110111";
		Trees_din <= x"ff650545";
		wait for Clk_period;
		Addr <=  "00000100111000";
		Trees_din <= x"1d004704";
		wait for Clk_period;
		Addr <=  "00000100111001";
		Trees_din <= x"00480545";
		wait for Clk_period;
		Addr <=  "00000100111010";
		Trees_din <= x"ffa30545";
		wait for Clk_period;
		Addr <=  "00000100111011";
		Trees_din <= x"1201910c";
		wait for Clk_period;
		Addr <=  "00000100111100";
		Trees_din <= x"04f70e04";
		wait for Clk_period;
		Addr <=  "00000100111101";
		Trees_din <= x"ffa70545";
		wait for Clk_period;
		Addr <=  "00000100111110";
		Trees_din <= x"08008104";
		wait for Clk_period;
		Addr <=  "00000100111111";
		Trees_din <= x"00910545";
		wait for Clk_period;
		Addr <=  "00000101000000";
		Trees_din <= x"000d0545";
		wait for Clk_period;
		Addr <=  "00000101000001";
		Trees_din <= x"ff880545";
		wait for Clk_period;
		Addr <=  "00000101000010";
		Trees_din <= x"06091b14";
		wait for Clk_period;
		Addr <=  "00000101000011";
		Trees_din <= x"11ff5e04";
		wait for Clk_period;
		Addr <=  "00000101000100";
		Trees_din <= x"ff9e0545";
		wait for Clk_period;
		Addr <=  "00000101000101";
		Trees_din <= x"0105950c";
		wait for Clk_period;
		Addr <=  "00000101000110";
		Trees_din <= x"0e00b204";
		wait for Clk_period;
		Addr <=  "00000101000111";
		Trees_din <= x"00940545";
		wait for Clk_period;
		Addr <=  "00000101001000";
		Trees_din <= x"14014e04";
		wait for Clk_period;
		Addr <=  "00000101001001";
		Trees_din <= x"ff900545";
		wait for Clk_period;
		Addr <=  "00000101001010";
		Trees_din <= x"00620545";
		wait for Clk_period;
		Addr <=  "00000101001011";
		Trees_din <= x"ffa80545";
		wait for Clk_period;
		Addr <=  "00000101001100";
		Trees_din <= x"0bfacb08";
		wait for Clk_period;
		Addr <=  "00000101001101";
		Trees_din <= x"06103104";
		wait for Clk_period;
		Addr <=  "00000101001110";
		Trees_din <= x"ffbf0545";
		wait for Clk_period;
		Addr <=  "00000101001111";
		Trees_din <= x"00770545";
		wait for Clk_period;
		Addr <=  "00000101010000";
		Trees_din <= x"00a20545";
		wait for Clk_period;
		Addr <=  "00000101010001";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00000101010010";
		Trees_din <= x"06023218";
		wait for Clk_period;
		Addr <=  "00000101010011";
		Trees_din <= x"06fee90c";
		wait for Clk_period;
		Addr <=  "00000101010100";
		Trees_din <= x"16040004";
		wait for Clk_period;
		Addr <=  "00000101010101";
		Trees_din <= x"ff6505bd";
		wait for Clk_period;
		Addr <=  "00000101010110";
		Trees_din <= x"13f87704";
		wait for Clk_period;
		Addr <=  "00000101010111";
		Trees_din <= x"004705bd";
		wait for Clk_period;
		Addr <=  "00000101011000";
		Trees_din <= x"ffa905bd";
		wait for Clk_period;
		Addr <=  "00000101011001";
		Trees_din <= x"0800e408";
		wait for Clk_period;
		Addr <=  "00000101011010";
		Trees_din <= x"08007804";
		wait for Clk_period;
		Addr <=  "00000101011011";
		Trees_din <= x"ffa805bd";
		wait for Clk_period;
		Addr <=  "00000101011100";
		Trees_din <= x"007105bd";
		wait for Clk_period;
		Addr <=  "00000101011101";
		Trees_din <= x"ff8c05bd";
		wait for Clk_period;
		Addr <=  "00000101011110";
		Trees_din <= x"06091b18";
		wait for Clk_period;
		Addr <=  "00000101011111";
		Trees_din <= x"1202000c";
		wait for Clk_period;
		Addr <=  "00000101100000";
		Trees_din <= x"04f9bb04";
		wait for Clk_period;
		Addr <=  "00000101100001";
		Trees_din <= x"ff8705bd";
		wait for Clk_period;
		Addr <=  "00000101100010";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00000101100011";
		Trees_din <= x"006505bd";
		wait for Clk_period;
		Addr <=  "00000101100100";
		Trees_din <= x"fff805bd";
		wait for Clk_period;
		Addr <=  "00000101100101";
		Trees_din <= x"09005604";
		wait for Clk_period;
		Addr <=  "00000101100110";
		Trees_din <= x"ffcc05bd";
		wait for Clk_period;
		Addr <=  "00000101100111";
		Trees_din <= x"19009104";
		wait for Clk_period;
		Addr <=  "00000101101000";
		Trees_din <= x"002505bd";
		wait for Clk_period;
		Addr <=  "00000101101001";
		Trees_din <= x"009205bd";
		wait for Clk_period;
		Addr <=  "00000101101010";
		Trees_din <= x"02009004";
		wait for Clk_period;
		Addr <=  "00000101101011";
		Trees_din <= x"009a05bd";
		wait for Clk_period;
		Addr <=  "00000101101100";
		Trees_din <= x"19008904";
		wait for Clk_period;
		Addr <=  "00000101101101";
		Trees_din <= x"005e05bd";
		wait for Clk_period;
		Addr <=  "00000101101110";
		Trees_din <= x"ffd005bd";
		wait for Clk_period;
		Addr <=  "00000101101111";
		Trees_din <= x"06023218";
		wait for Clk_period;
		Addr <=  "00000101110000";
		Trees_din <= x"06fee90c";
		wait for Clk_period;
		Addr <=  "00000101110001";
		Trees_din <= x"1703fd04";
		wait for Clk_period;
		Addr <=  "00000101110010";
		Trees_din <= x"ff660631";
		wait for Clk_period;
		Addr <=  "00000101110011";
		Trees_din <= x"0efe8f04";
		wait for Clk_period;
		Addr <=  "00000101110100";
		Trees_din <= x"00460631";
		wait for Clk_period;
		Addr <=  "00000101110101";
		Trees_din <= x"ffad0631";
		wait for Clk_period;
		Addr <=  "00000101110110";
		Trees_din <= x"0800e408";
		wait for Clk_period;
		Addr <=  "00000101110111";
		Trees_din <= x"08007804";
		wait for Clk_period;
		Addr <=  "00000101111000";
		Trees_din <= x"ffae0631";
		wait for Clk_period;
		Addr <=  "00000101111001";
		Trees_din <= x"00660631";
		wait for Clk_period;
		Addr <=  "00000101111010";
		Trees_din <= x"ff900631";
		wait for Clk_period;
		Addr <=  "00000101111011";
		Trees_din <= x"06091b18";
		wait for Clk_period;
		Addr <=  "00000101111100";
		Trees_din <= x"12024310";
		wait for Clk_period;
		Addr <=  "00000101111101";
		Trees_din <= x"04f9bb08";
		wait for Clk_period;
		Addr <=  "00000101111110";
		Trees_din <= x"05f8f704";
		wait for Clk_period;
		Addr <=  "00000101111111";
		Trees_din <= x"fffc0631";
		wait for Clk_period;
		Addr <=  "00000110000000";
		Trees_din <= x"ff930631";
		wait for Clk_period;
		Addr <=  "00000110000001";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "00000110000010";
		Trees_din <= x"00440631";
		wait for Clk_period;
		Addr <=  "00000110000011";
		Trees_din <= x"fff40631";
		wait for Clk_period;
		Addr <=  "00000110000100";
		Trees_din <= x"09005604";
		wait for Clk_period;
		Addr <=  "00000110000101";
		Trees_din <= x"00030631";
		wait for Clk_period;
		Addr <=  "00000110000110";
		Trees_din <= x"00720631";
		wait for Clk_period;
		Addr <=  "00000110000111";
		Trees_din <= x"0bfacb08";
		wait for Clk_period;
		Addr <=  "00000110001000";
		Trees_din <= x"06103104";
		wait for Clk_period;
		Addr <=  "00000110001001";
		Trees_din <= x"ffbd0631";
		wait for Clk_period;
		Addr <=  "00000110001010";
		Trees_din <= x"00680631";
		wait for Clk_period;
		Addr <=  "00000110001011";
		Trees_din <= x"009a0631";
		wait for Clk_period;
		Addr <=  "00000110001100";
		Trees_din <= x"06ffc30c";
		wait for Clk_period;
		Addr <=  "00000110001101";
		Trees_din <= x"16040008";
		wait for Clk_period;
		Addr <=  "00000110001110";
		Trees_din <= x"06fee904";
		wait for Clk_period;
		Addr <=  "00000110001111";
		Trees_din <= x"ff66068d";
		wait for Clk_period;
		Addr <=  "00000110010000";
		Trees_din <= x"ffe1068d";
		wait for Clk_period;
		Addr <=  "00000110010001";
		Trees_din <= x"fffd068d";
		wait for Clk_period;
		Addr <=  "00000110010010";
		Trees_din <= x"06091b18";
		wait for Clk_period;
		Addr <=  "00000110010011";
		Trees_din <= x"04f4a204";
		wait for Clk_period;
		Addr <=  "00000110010100";
		Trees_din <= x"ff99068d";
		wait for Clk_period;
		Addr <=  "00000110010101";
		Trees_din <= x"0f010808";
		wait for Clk_period;
		Addr <=  "00000110010110";
		Trees_din <= x"1603d904";
		wait for Clk_period;
		Addr <=  "00000110010111";
		Trees_din <= x"ff95068d";
		wait for Clk_period;
		Addr <=  "00000110011000";
		Trees_din <= x"0026068d";
		wait for Clk_period;
		Addr <=  "00000110011001";
		Trees_din <= x"07005908";
		wait for Clk_period;
		Addr <=  "00000110011010";
		Trees_din <= x"12010f04";
		wait for Clk_period;
		Addr <=  "00000110011011";
		Trees_din <= x"0001068d";
		wait for Clk_period;
		Addr <=  "00000110011100";
		Trees_din <= x"008e068d";
		wait for Clk_period;
		Addr <=  "00000110011101";
		Trees_din <= x"ffe3068d";
		wait for Clk_period;
		Addr <=  "00000110011110";
		Trees_din <= x"0bfacb08";
		wait for Clk_period;
		Addr <=  "00000110011111";
		Trees_din <= x"06103104";
		wait for Clk_period;
		Addr <=  "00000110100000";
		Trees_din <= x"ffc0068d";
		wait for Clk_period;
		Addr <=  "00000110100001";
		Trees_din <= x"0060068d";
		wait for Clk_period;
		Addr <=  "00000110100010";
		Trees_din <= x"0095068d";
		wait for Clk_period;
		Addr <=  "00000110100011";
		Trees_din <= x"06fee908";
		wait for Clk_period;
		Addr <=  "00000110100100";
		Trees_din <= x"1703fd04";
		wait for Clk_period;
		Addr <=  "00000110100101";
		Trees_din <= x"ff6706e1";
		wait for Clk_period;
		Addr <=  "00000110100110";
		Trees_din <= x"000406e1";
		wait for Clk_period;
		Addr <=  "00000110100111";
		Trees_din <= x"06091b18";
		wait for Clk_period;
		Addr <=  "00000110101000";
		Trees_din <= x"01060b14";
		wait for Clk_period;
		Addr <=  "00000110101001";
		Trees_din <= x"0f00ff08";
		wait for Clk_period;
		Addr <=  "00000110101010";
		Trees_din <= x"0f000f04";
		wait for Clk_period;
		Addr <=  "00000110101011";
		Trees_din <= x"001806e1";
		wait for Clk_period;
		Addr <=  "00000110101100";
		Trees_din <= x"ffa406e1";
		wait for Clk_period;
		Addr <=  "00000110101101";
		Trees_din <= x"1b003104";
		wait for Clk_period;
		Addr <=  "00000110101110";
		Trees_din <= x"ffcf06e1";
		wait for Clk_period;
		Addr <=  "00000110101111";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00000110110000";
		Trees_din <= x"007f06e1";
		wait for Clk_period;
		Addr <=  "00000110110001";
		Trees_din <= x"ffe906e1";
		wait for Clk_period;
		Addr <=  "00000110110010";
		Trees_din <= x"ff9a06e1";
		wait for Clk_period;
		Addr <=  "00000110110011";
		Trees_din <= x"0bfacb08";
		wait for Clk_period;
		Addr <=  "00000110110100";
		Trees_din <= x"06103104";
		wait for Clk_period;
		Addr <=  "00000110110101";
		Trees_din <= x"ffc406e1";
		wait for Clk_period;
		Addr <=  "00000110110110";
		Trees_din <= x"005a06e1";
		wait for Clk_period;
		Addr <=  "00000110110111";
		Trees_din <= x"009106e1";
		wait for Clk_period;
		Addr <=  "00000110111000";
		Trees_din <= x"06ffc30c";
		wait for Clk_period;
		Addr <=  "00000110111001";
		Trees_din <= x"16040008";
		wait for Clk_period;
		Addr <=  "00000110111010";
		Trees_din <= x"06fee904";
		wait for Clk_period;
		Addr <=  "00000110111011";
		Trees_din <= x"ff67073d";
		wait for Clk_period;
		Addr <=  "00000110111100";
		Trees_din <= x"ffe2073d";
		wait for Clk_period;
		Addr <=  "00000110111101";
		Trees_din <= x"0007073d";
		wait for Clk_period;
		Addr <=  "00000110111110";
		Trees_din <= x"06091b18";
		wait for Clk_period;
		Addr <=  "00000110111111";
		Trees_din <= x"04f9a010";
		wait for Clk_period;
		Addr <=  "00000111000000";
		Trees_din <= x"16006908";
		wait for Clk_period;
		Addr <=  "00000111000001";
		Trees_din <= x"07005704";
		wait for Clk_period;
		Addr <=  "00000111000010";
		Trees_din <= x"0064073d";
		wait for Clk_period;
		Addr <=  "00000111000011";
		Trees_din <= x"fff2073d";
		wait for Clk_period;
		Addr <=  "00000111000100";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00000111000101";
		Trees_din <= x"ff89073d";
		wait for Clk_period;
		Addr <=  "00000111000110";
		Trees_din <= x"ffed073d";
		wait for Clk_period;
		Addr <=  "00000111000111";
		Trees_din <= x"00fd2504";
		wait for Clk_period;
		Addr <=  "00000111001000";
		Trees_din <= x"fff7073d";
		wait for Clk_period;
		Addr <=  "00000111001001";
		Trees_din <= x"0061073d";
		wait for Clk_period;
		Addr <=  "00000111001010";
		Trees_din <= x"0bfacb08";
		wait for Clk_period;
		Addr <=  "00000111001011";
		Trees_din <= x"06103104";
		wait for Clk_period;
		Addr <=  "00000111001100";
		Trees_din <= x"ffc8073d";
		wait for Clk_period;
		Addr <=  "00000111001101";
		Trees_din <= x"0053073d";
		wait for Clk_period;
		Addr <=  "00000111001110";
		Trees_din <= x"008c073d";
		wait for Clk_period;
		Addr <=  "00000111001111";
		Trees_din <= x"06ffc30c";
		wait for Clk_period;
		Addr <=  "00000111010000";
		Trees_din <= x"1703fd08";
		wait for Clk_period;
		Addr <=  "00000111010001";
		Trees_din <= x"06fee904";
		wait for Clk_period;
		Addr <=  "00000111010010";
		Trees_din <= x"ff680791";
		wait for Clk_period;
		Addr <=  "00000111010011";
		Trees_din <= x"ffe30791";
		wait for Clk_period;
		Addr <=  "00000111010100";
		Trees_din <= x"000d0791";
		wait for Clk_period;
		Addr <=  "00000111010101";
		Trees_din <= x"06091b18";
		wait for Clk_period;
		Addr <=  "00000111010110";
		Trees_din <= x"01060b14";
		wait for Clk_period;
		Addr <=  "00000111010111";
		Trees_din <= x"0c028d0c";
		wait for Clk_period;
		Addr <=  "00000111011000";
		Trees_din <= x"01034108";
		wait for Clk_period;
		Addr <=  "00000111011001";
		Trees_din <= x"1900a004";
		wait for Clk_period;
		Addr <=  "00000111011010";
		Trees_din <= x"ffa20791";
		wait for Clk_period;
		Addr <=  "00000111011011";
		Trees_din <= x"00060791";
		wait for Clk_period;
		Addr <=  "00000111011100";
		Trees_din <= x"00530791";
		wait for Clk_period;
		Addr <=  "00000111011101";
		Trees_din <= x"05fbfd04";
		wait for Clk_period;
		Addr <=  "00000111011110";
		Trees_din <= x"00220791";
		wait for Clk_period;
		Addr <=  "00000111011111";
		Trees_din <= x"006f0791";
		wait for Clk_period;
		Addr <=  "00000111100000";
		Trees_din <= x"ffa60791";
		wait for Clk_period;
		Addr <=  "00000111100001";
		Trees_din <= x"02009004";
		wait for Clk_period;
		Addr <=  "00000111100010";
		Trees_din <= x"00820791";
		wait for Clk_period;
		Addr <=  "00000111100011";
		Trees_din <= x"00030791";
		wait for Clk_period;
		Addr <=  "00000111100100";
		Trees_din <= x"06fee908";
		wait for Clk_period;
		Addr <=  "00000111100101";
		Trees_din <= x"16040004";
		wait for Clk_period;
		Addr <=  "00000111100110";
		Trees_din <= x"ff6907e5";
		wait for Clk_period;
		Addr <=  "00000111100111";
		Trees_din <= x"000f07e5";
		wait for Clk_period;
		Addr <=  "00000111101000";
		Trees_din <= x"00046418";
		wait for Clk_period;
		Addr <=  "00000111101001";
		Trees_din <= x"07005004";
		wait for Clk_period;
		Addr <=  "00000111101010";
		Trees_din <= x"ffd607e5";
		wait for Clk_period;
		Addr <=  "00000111101011";
		Trees_din <= x"06091b10";
		wait for Clk_period;
		Addr <=  "00000111101100";
		Trees_din <= x"07005908";
		wait for Clk_period;
		Addr <=  "00000111101101";
		Trees_din <= x"0f00fb04";
		wait for Clk_period;
		Addr <=  "00000111101110";
		Trees_din <= x"fff807e5";
		wait for Clk_period;
		Addr <=  "00000111101111";
		Trees_din <= x"006807e5";
		wait for Clk_period;
		Addr <=  "00000111110000";
		Trees_din <= x"1c003904";
		wait for Clk_period;
		Addr <=  "00000111110001";
		Trees_din <= x"001907e5";
		wait for Clk_period;
		Addr <=  "00000111110010";
		Trees_din <= x"ffc107e5";
		wait for Clk_period;
		Addr <=  "00000111110011";
		Trees_din <= x"008407e5";
		wait for Clk_period;
		Addr <=  "00000111110100";
		Trees_din <= x"02ffb908";
		wait for Clk_period;
		Addr <=  "00000111110101";
		Trees_din <= x"09005804";
		wait for Clk_period;
		Addr <=  "00000111110110";
		Trees_din <= x"ffea07e5";
		wait for Clk_period;
		Addr <=  "00000111110111";
		Trees_din <= x"004a07e5";
		wait for Clk_period;
		Addr <=  "00000111111000";
		Trees_din <= x"ff8f07e5";
		wait for Clk_period;
		Addr <=  "00000111111001";
		Trees_din <= x"06fee908";
		wait for Clk_period;
		Addr <=  "00000111111010";
		Trees_din <= x"1703fd04";
		wait for Clk_period;
		Addr <=  "00000111111011";
		Trees_din <= x"ff6a0839";
		wait for Clk_period;
		Addr <=  "00000111111100";
		Trees_din <= x"00150839";
		wait for Clk_period;
		Addr <=  "00000111111101";
		Trees_din <= x"00046418";
		wait for Clk_period;
		Addr <=  "00000111111110";
		Trees_din <= x"06091b14";
		wait for Clk_period;
		Addr <=  "00000111111111";
		Trees_din <= x"14012e08";
		wait for Clk_period;
		Addr <=  "00001000000000";
		Trees_din <= x"13fdce04";
		wait for Clk_period;
		Addr <=  "00001000000001";
		Trees_din <= x"00110839";
		wait for Clk_period;
		Addr <=  "00001000000010";
		Trees_din <= x"ffa60839";
		wait for Clk_period;
		Addr <=  "00001000000011";
		Trees_din <= x"08017508";
		wait for Clk_period;
		Addr <=  "00001000000100";
		Trees_din <= x"07005704";
		wait for Clk_period;
		Addr <=  "00001000000101";
		Trees_din <= x"00710839";
		wait for Clk_period;
		Addr <=  "00001000000110";
		Trees_din <= x"00140839";
		wait for Clk_period;
		Addr <=  "00001000000111";
		Trees_din <= x"fff10839";
		wait for Clk_period;
		Addr <=  "00001000001000";
		Trees_din <= x"00750839";
		wait for Clk_period;
		Addr <=  "00001000001001";
		Trees_din <= x"02ffb908";
		wait for Clk_period;
		Addr <=  "00001000001010";
		Trees_din <= x"09005804";
		wait for Clk_period;
		Addr <=  "00001000001011";
		Trees_din <= x"ffeb0839";
		wait for Clk_period;
		Addr <=  "00001000001100";
		Trees_din <= x"00460839";
		wait for Clk_period;
		Addr <=  "00001000001101";
		Trees_din <= x"ff940839";
		wait for Clk_period;
		Addr <=  "00001000001110";
		Trees_din <= x"06ffc30c";
		wait for Clk_period;
		Addr <=  "00001000001111";
		Trees_din <= x"16040008";
		wait for Clk_period;
		Addr <=  "00001000010000";
		Trees_din <= x"06fee904";
		wait for Clk_period;
		Addr <=  "00001000010001";
		Trees_din <= x"ff6a0885";
		wait for Clk_period;
		Addr <=  "00001000010010";
		Trees_din <= x"ffe40885";
		wait for Clk_period;
		Addr <=  "00001000010011";
		Trees_din <= x"00180885";
		wait for Clk_period;
		Addr <=  "00001000010100";
		Trees_din <= x"01060b14";
		wait for Clk_period;
		Addr <=  "00001000010101";
		Trees_din <= x"00068110";
		wait for Clk_period;
		Addr <=  "00001000010110";
		Trees_din <= x"06091b0c";
		wait for Clk_period;
		Addr <=  "00001000010111";
		Trees_din <= x"14014604";
		wait for Clk_period;
		Addr <=  "00001000011000";
		Trees_din <= x"ffd90885";
		wait for Clk_period;
		Addr <=  "00001000011001";
		Trees_din <= x"00fd2504";
		wait for Clk_period;
		Addr <=  "00001000011010";
		Trees_din <= x"fffc0885";
		wait for Clk_period;
		Addr <=  "00001000011011";
		Trees_din <= x"00690885";
		wait for Clk_period;
		Addr <=  "00001000011100";
		Trees_din <= x"007b0885";
		wait for Clk_period;
		Addr <=  "00001000011101";
		Trees_din <= x"ffe50885";
		wait for Clk_period;
		Addr <=  "00001000011110";
		Trees_din <= x"16026f04";
		wait for Clk_period;
		Addr <=  "00001000011111";
		Trees_din <= x"fffe0885";
		wait for Clk_period;
		Addr <=  "00001000100000";
		Trees_din <= x"ffb70885";
		wait for Clk_period;
		Addr <=  "00001000100001";
		Trees_din <= x"06fee908";
		wait for Clk_period;
		Addr <=  "00001000100010";
		Trees_din <= x"1703fd04";
		wait for Clk_period;
		Addr <=  "00001000100011";
		Trees_din <= x"ff6b08c9";
		wait for Clk_period;
		Addr <=  "00001000100100";
		Trees_din <= x"001908c9";
		wait for Clk_period;
		Addr <=  "00001000100101";
		Trees_din <= x"02002410";
		wait for Clk_period;
		Addr <=  "00001000100110";
		Trees_din <= x"05fdb60c";
		wait for Clk_period;
		Addr <=  "00001000100111";
		Trees_din <= x"0d031708";
		wait for Clk_period;
		Addr <=  "00001000101000";
		Trees_din <= x"1c003b04";
		wait for Clk_period;
		Addr <=  "00001000101001";
		Trees_din <= x"007108c9";
		wait for Clk_period;
		Addr <=  "00001000101010";
		Trees_din <= x"001c08c9";
		wait for Clk_period;
		Addr <=  "00001000101011";
		Trees_din <= x"fff908c9";
		wait for Clk_period;
		Addr <=  "00001000101100";
		Trees_din <= x"ffde08c9";
		wait for Clk_period;
		Addr <=  "00001000101101";
		Trees_din <= x"0002d308";
		wait for Clk_period;
		Addr <=  "00001000101110";
		Trees_din <= x"00fe2904";
		wait for Clk_period;
		Addr <=  "00001000101111";
		Trees_din <= x"ffda08c9";
		wait for Clk_period;
		Addr <=  "00001000110000";
		Trees_din <= x"004808c9";
		wait for Clk_period;
		Addr <=  "00001000110001";
		Trees_din <= x"ff9908c9";
		wait for Clk_period;
		Addr <=  "00001000110010";
		Trees_din <= x"06f9ca04";
		wait for Clk_period;
		Addr <=  "00001000110011";
		Trees_din <= x"ff6d0915";
		wait for Clk_period;
		Addr <=  "00001000110100";
		Trees_din <= x"0003e518";
		wait for Clk_period;
		Addr <=  "00001000110101";
		Trees_din <= x"13f96908";
		wait for Clk_period;
		Addr <=  "00001000110110";
		Trees_din <= x"02fe8304";
		wait for Clk_period;
		Addr <=  "00001000110111";
		Trees_din <= x"00a00915";
		wait for Clk_period;
		Addr <=  "00001000111000";
		Trees_din <= x"000f0915";
		wait for Clk_period;
		Addr <=  "00001000111001";
		Trees_din <= x"06054008";
		wait for Clk_period;
		Addr <=  "00001000111010";
		Trees_din <= x"1e006e04";
		wait for Clk_period;
		Addr <=  "00001000111011";
		Trees_din <= x"ffa40915";
		wait for Clk_period;
		Addr <=  "00001000111100";
		Trees_din <= x"000c0915";
		wait for Clk_period;
		Addr <=  "00001000111101";
		Trees_din <= x"1701d504";
		wait for Clk_period;
		Addr <=  "00001000111110";
		Trees_din <= x"00630915";
		wait for Clk_period;
		Addr <=  "00001000111111";
		Trees_din <= x"fff10915";
		wait for Clk_period;
		Addr <=  "00001001000000";
		Trees_din <= x"06023204";
		wait for Clk_period;
		Addr <=  "00001001000001";
		Trees_din <= x"ff8a0915";
		wait for Clk_period;
		Addr <=  "00001001000010";
		Trees_din <= x"11024c04";
		wait for Clk_period;
		Addr <=  "00001001000011";
		Trees_din <= x"ffd00915";
		wait for Clk_period;
		Addr <=  "00001001000100";
		Trees_din <= x"00370915";
		wait for Clk_period;
		Addr <=  "00001001000101";
		Trees_din <= x"06f9ca04";
		wait for Clk_period;
		Addr <=  "00001001000110";
		Trees_din <= x"ff6e0961";
		wait for Clk_period;
		Addr <=  "00001001000111";
		Trees_din <= x"0003e518";
		wait for Clk_period;
		Addr <=  "00001001001000";
		Trees_din <= x"18004610";
		wait for Clk_period;
		Addr <=  "00001001001001";
		Trees_din <= x"06054008";
		wait for Clk_period;
		Addr <=  "00001001001010";
		Trees_din <= x"12fecd04";
		wait for Clk_period;
		Addr <=  "00001001001011";
		Trees_din <= x"00180961";
		wait for Clk_period;
		Addr <=  "00001001001100";
		Trees_din <= x"ffa40961";
		wait for Clk_period;
		Addr <=  "00001001001101";
		Trees_din <= x"1701d504";
		wait for Clk_period;
		Addr <=  "00001001001110";
		Trees_din <= x"00590961";
		wait for Clk_period;
		Addr <=  "00001001001111";
		Trees_din <= x"fff90961";
		wait for Clk_period;
		Addr <=  "00001001010000";
		Trees_din <= x"1e007804";
		wait for Clk_period;
		Addr <=  "00001001010001";
		Trees_din <= x"009b0961";
		wait for Clk_period;
		Addr <=  "00001001010010";
		Trees_din <= x"001a0961";
		wait for Clk_period;
		Addr <=  "00001001010011";
		Trees_din <= x"02ffb908";
		wait for Clk_period;
		Addr <=  "00001001010100";
		Trees_din <= x"09005804";
		wait for Clk_period;
		Addr <=  "00001001010101";
		Trees_din <= x"ffd80961";
		wait for Clk_period;
		Addr <=  "00001001010110";
		Trees_din <= x"00350961";
		wait for Clk_period;
		Addr <=  "00001001010111";
		Trees_din <= x"ff8c0961";
		wait for Clk_period;
		Addr <=  "00001001011000";
		Trees_din <= x"06f9ca04";
		wait for Clk_period;
		Addr <=  "00001001011001";
		Trees_din <= x"ff6f09a5";
		wait for Clk_period;
		Addr <=  "00001001011010";
		Trees_din <= x"13f9690c";
		wait for Clk_period;
		Addr <=  "00001001011011";
		Trees_din <= x"02ffb908";
		wait for Clk_period;
		Addr <=  "00001001011100";
		Trees_din <= x"0d003004";
		wait for Clk_period;
		Addr <=  "00001001011101";
		Trees_din <= x"009809a5";
		wait for Clk_period;
		Addr <=  "00001001011110";
		Trees_din <= x"002509a5";
		wait for Clk_period;
		Addr <=  "00001001011111";
		Trees_din <= x"fff909a5";
		wait for Clk_period;
		Addr <=  "00001001100000";
		Trees_din <= x"06054008";
		wait for Clk_period;
		Addr <=  "00001001100001";
		Trees_din <= x"0afae404";
		wait for Clk_period;
		Addr <=  "00001001100010";
		Trees_din <= x"ffe409a5";
		wait for Clk_period;
		Addr <=  "00001001100011";
		Trees_din <= x"ff8c09a5";
		wait for Clk_period;
		Addr <=  "00001001100100";
		Trees_din <= x"14014e04";
		wait for Clk_period;
		Addr <=  "00001001100101";
		Trees_din <= x"ffe609a5";
		wait for Clk_period;
		Addr <=  "00001001100110";
		Trees_din <= x"12018b04";
		wait for Clk_period;
		Addr <=  "00001001100111";
		Trees_din <= x"000209a5";
		wait for Clk_period;
		Addr <=  "00001001101000";
		Trees_din <= x"006809a5";
		wait for Clk_period;
		Addr <=  "00001001101001";
		Trees_din <= x"06f9ca04";
		wait for Clk_period;
		Addr <=  "00001001101010";
		Trees_din <= x"ff7109e9";
		wait for Clk_period;
		Addr <=  "00001001101011";
		Trees_din <= x"0003e514";
		wait for Clk_period;
		Addr <=  "00001001101100";
		Trees_din <= x"14002604";
		wait for Clk_period;
		Addr <=  "00001001101101";
		Trees_din <= x"008709e9";
		wait for Clk_period;
		Addr <=  "00001001101110";
		Trees_din <= x"06091b0c";
		wait for Clk_period;
		Addr <=  "00001001101111";
		Trees_din <= x"0f00ff04";
		wait for Clk_period;
		Addr <=  "00001001110000";
		Trees_din <= x"ffb209e9";
		wait for Clk_period;
		Addr <=  "00001001110001";
		Trees_din <= x"07005904";
		wait for Clk_period;
		Addr <=  "00001001110010";
		Trees_din <= x"004509e9";
		wait for Clk_period;
		Addr <=  "00001001110011";
		Trees_din <= x"ffdd09e9";
		wait for Clk_period;
		Addr <=  "00001001110100";
		Trees_din <= x"005609e9";
		wait for Clk_period;
		Addr <=  "00001001110101";
		Trees_din <= x"02ffb908";
		wait for Clk_period;
		Addr <=  "00001001110110";
		Trees_din <= x"04f73904";
		wait for Clk_period;
		Addr <=  "00001001110111";
		Trees_din <= x"003309e9";
		wait for Clk_period;
		Addr <=  "00001001111000";
		Trees_din <= x"ffd809e9";
		wait for Clk_period;
		Addr <=  "00001001111001";
		Trees_din <= x"ff9309e9";
		wait for Clk_period;
		Addr <=  "00001001111010";
		Trees_din <= x"06f9ca04";
		wait for Clk_period;
		Addr <=  "00001001111011";
		Trees_din <= x"ff730a25";
		wait for Clk_period;
		Addr <=  "00001001111100";
		Trees_din <= x"13f96908";
		wait for Clk_period;
		Addr <=  "00001001111101";
		Trees_din <= x"02ffb904";
		wait for Clk_period;
		Addr <=  "00001001111110";
		Trees_din <= x"00770a25";
		wait for Clk_period;
		Addr <=  "00001001111111";
		Trees_din <= x"fffc0a25";
		wait for Clk_period;
		Addr <=  "00001010000000";
		Trees_din <= x"06054008";
		wait for Clk_period;
		Addr <=  "00001010000001";
		Trees_din <= x"18004604";
		wait for Clk_period;
		Addr <=  "00001010000010";
		Trees_din <= x"ff910a25";
		wait for Clk_period;
		Addr <=  "00001010000011";
		Trees_din <= x"ffea0a25";
		wait for Clk_period;
		Addr <=  "00001010000100";
		Trees_din <= x"04f47104";
		wait for Clk_period;
		Addr <=  "00001010000101";
		Trees_din <= x"ffdb0a25";
		wait for Clk_period;
		Addr <=  "00001010000110";
		Trees_din <= x"11023604";
		wait for Clk_period;
		Addr <=  "00001010000111";
		Trees_din <= x"ffff0a25";
		wait for Clk_period;
		Addr <=  "00001010001000";
		Trees_din <= x"00550a25";
		wait for Clk_period;
		Addr <=  "00001010001001";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "00001010001010";
		Trees_din <= x"06f9ca04";
		wait for Clk_period;
		Addr <=  "00001010001011";
		Trees_din <= x"ff750a65";
		wait for Clk_period;
		Addr <=  "00001010001100";
		Trees_din <= x"0003e514";
		wait for Clk_period;
		Addr <=  "00001010001101";
		Trees_din <= x"0a020f0c";
		wait for Clk_period;
		Addr <=  "00001010001110";
		Trees_din <= x"06091b08";
		wait for Clk_period;
		Addr <=  "00001010001111";
		Trees_din <= x"01039c04";
		wait for Clk_period;
		Addr <=  "00001010010000";
		Trees_din <= x"ffbe0a65";
		wait for Clk_period;
		Addr <=  "00001010010001";
		Trees_din <= x"00260a65";
		wait for Clk_period;
		Addr <=  "00001010010010";
		Trees_din <= x"003d0a65";
		wait for Clk_period;
		Addr <=  "00001010010011";
		Trees_din <= x"0a027604";
		wait for Clk_period;
		Addr <=  "00001010010100";
		Trees_din <= x"00880a65";
		wait for Clk_period;
		Addr <=  "00001010010101";
		Trees_din <= x"00170a65";
		wait for Clk_period;
		Addr <=  "00001010010110";
		Trees_din <= x"06023204";
		wait for Clk_period;
		Addr <=  "00001010010111";
		Trees_din <= x"ff9b0a65";
		wait for Clk_period;
		Addr <=  "00001010011000";
		Trees_din <= x"00090a65";
		wait for Clk_period;
		Addr <=  "00001010011001";
		Trees_din <= x"06f9ca04";
		wait for Clk_period;
		Addr <=  "00001010011010";
		Trees_din <= x"ff770aa1";
		wait for Clk_period;
		Addr <=  "00001010011011";
		Trees_din <= x"00068114";
		wait for Clk_period;
		Addr <=  "00001010011100";
		Trees_din <= x"01070110";
		wait for Clk_period;
		Addr <=  "00001010011101";
		Trees_din <= x"05fdb60c";
		wait for Clk_period;
		Addr <=  "00001010011110";
		Trees_din <= x"1b003504";
		wait for Clk_period;
		Addr <=  "00001010011111";
		Trees_din <= x"ffff0aa1";
		wait for Clk_period;
		Addr <=  "00001010100000";
		Trees_din <= x"1a00b404";
		wait for Clk_period;
		Addr <=  "00001010100001";
		Trees_din <= x"001e0aa1";
		wait for Clk_period;
		Addr <=  "00001010100010";
		Trees_din <= x"00760aa1";
		wait for Clk_period;
		Addr <=  "00001010100011";
		Trees_din <= x"fff30aa1";
		wait for Clk_period;
		Addr <=  "00001010100100";
		Trees_din <= x"ffc90aa1";
		wait for Clk_period;
		Addr <=  "00001010100101";
		Trees_din <= x"12027d04";
		wait for Clk_period;
		Addr <=  "00001010100110";
		Trees_din <= x"ffa40aa1";
		wait for Clk_period;
		Addr <=  "00001010100111";
		Trees_din <= x"fffe0aa1";
		wait for Clk_period;
		Addr <=  "00001010101000";
		Trees_din <= x"06f9ca04";
		wait for Clk_period;
		Addr <=  "00001010101001";
		Trees_din <= x"ff790add";
		wait for Clk_period;
		Addr <=  "00001010101010";
		Trees_din <= x"13f96908";
		wait for Clk_period;
		Addr <=  "00001010101011";
		Trees_din <= x"02ffb904";
		wait for Clk_period;
		Addr <=  "00001010101100";
		Trees_din <= x"00670add";
		wait for Clk_period;
		Addr <=  "00001010101101";
		Trees_din <= x"fffb0add";
		wait for Clk_period;
		Addr <=  "00001010101110";
		Trees_din <= x"06054008";
		wait for Clk_period;
		Addr <=  "00001010101111";
		Trees_din <= x"0afae404";
		wait for Clk_period;
		Addr <=  "00001010110000";
		Trees_din <= x"ffee0add";
		wait for Clk_period;
		Addr <=  "00001010110001";
		Trees_din <= x"ff990add";
		wait for Clk_period;
		Addr <=  "00001010110010";
		Trees_din <= x"04f47104";
		wait for Clk_period;
		Addr <=  "00001010110011";
		Trees_din <= x"ffdf0add";
		wait for Clk_period;
		Addr <=  "00001010110100";
		Trees_din <= x"12019704";
		wait for Clk_period;
		Addr <=  "00001010110101";
		Trees_din <= x"00090add";
		wait for Clk_period;
		Addr <=  "00001010110110";
		Trees_din <= x"00460add";
		wait for Clk_period;
		Addr <=  "00001010110111";
		Trees_din <= x"06f9ca04";
		wait for Clk_period;
		Addr <=  "00001010111000";
		Trees_din <= x"ff7c0b19";
		wait for Clk_period;
		Addr <=  "00001010111001";
		Trees_din <= x"0004a114";
		wait for Clk_period;
		Addr <=  "00001010111010";
		Trees_din <= x"1800460c";
		wait for Clk_period;
		Addr <=  "00001010111011";
		Trees_din <= x"06091b08";
		wait for Clk_period;
		Addr <=  "00001010111100";
		Trees_din <= x"0d02f204";
		wait for Clk_period;
		Addr <=  "00001010111101";
		Trees_din <= x"ffc20b19";
		wait for Clk_period;
		Addr <=  "00001010111110";
		Trees_din <= x"00110b19";
		wait for Clk_period;
		Addr <=  "00001010111111";
		Trees_din <= x"003a0b19";
		wait for Clk_period;
		Addr <=  "00001011000000";
		Trees_din <= x"1e007804";
		wait for Clk_period;
		Addr <=  "00001011000001";
		Trees_din <= x"006e0b19";
		wait for Clk_period;
		Addr <=  "00001011000010";
		Trees_din <= x"000c0b19";
		wait for Clk_period;
		Addr <=  "00001011000011";
		Trees_din <= x"02ffb904";
		wait for Clk_period;
		Addr <=  "00001011000100";
		Trees_din <= x"00040b19";
		wait for Clk_period;
		Addr <=  "00001011000101";
		Trees_din <= x"ffa20b19";
		wait for Clk_period;
		Addr <=  "00001011000110";
		Trees_din <= x"06f9ca04";
		wait for Clk_period;
		Addr <=  "00001011000111";
		Trees_din <= x"ff7f0b55";
		wait for Clk_period;
		Addr <=  "00001011001000";
		Trees_din <= x"00068114";
		wait for Clk_period;
		Addr <=  "00001011001001";
		Trees_din <= x"01070110";
		wait for Clk_period;
		Addr <=  "00001011001010";
		Trees_din <= x"05fdb60c";
		wait for Clk_period;
		Addr <=  "00001011001011";
		Trees_din <= x"0200e808";
		wait for Clk_period;
		Addr <=  "00001011001100";
		Trees_din <= x"01fe6a04";
		wait for Clk_period;
		Addr <=  "00001011001101";
		Trees_din <= x"00050b55";
		wait for Clk_period;
		Addr <=  "00001011001110";
		Trees_din <= x"00700b55";
		wait for Clk_period;
		Addr <=  "00001011001111";
		Trees_din <= x"ffff0b55";
		wait for Clk_period;
		Addr <=  "00001011010000";
		Trees_din <= x"fff30b55";
		wait for Clk_period;
		Addr <=  "00001011010001";
		Trees_din <= x"ffcd0b55";
		wait for Clk_period;
		Addr <=  "00001011010010";
		Trees_din <= x"03f89804";
		wait for Clk_period;
		Addr <=  "00001011010011";
		Trees_din <= x"fff30b55";
		wait for Clk_period;
		Addr <=  "00001011010100";
		Trees_din <= x"ffaf0b55";
		wait for Clk_period;
		Addr <=  "00001011010101";
		Trees_din <= x"06f9ca04";
		wait for Clk_period;
		Addr <=  "00001011010110";
		Trees_din <= x"ff820b91";
		wait for Clk_period;
		Addr <=  "00001011010111";
		Trees_din <= x"13f96908";
		wait for Clk_period;
		Addr <=  "00001011011000";
		Trees_din <= x"02fe0104";
		wait for Clk_period;
		Addr <=  "00001011011001";
		Trees_din <= x"00600b91";
		wait for Clk_period;
		Addr <=  "00001011011010";
		Trees_din <= x"00030b91";
		wait for Clk_period;
		Addr <=  "00001011011011";
		Trees_din <= x"06054008";
		wait for Clk_period;
		Addr <=  "00001011011100";
		Trees_din <= x"1e007004";
		wait for Clk_period;
		Addr <=  "00001011011101";
		Trees_din <= x"ffa10b91";
		wait for Clk_period;
		Addr <=  "00001011011110";
		Trees_din <= x"ffe70b91";
		wait for Clk_period;
		Addr <=  "00001011011111";
		Trees_din <= x"14014e04";
		wait for Clk_period;
		Addr <=  "00001011100000";
		Trees_din <= x"ffe60b91";
		wait for Clk_period;
		Addr <=  "00001011100001";
		Trees_din <= x"10fdbe04";
		wait for Clk_period;
		Addr <=  "00001011100010";
		Trees_din <= x"00440b91";
		wait for Clk_period;
		Addr <=  "00001011100011";
		Trees_din <= x"00110b91";
		wait for Clk_period;
		Addr <=  "00001011100100";
		Trees_din <= x"06f9ca04";
		wait for Clk_period;
		Addr <=  "00001011100101";
		Trees_din <= x"ff850bc5";
		wait for Clk_period;
		Addr <=  "00001011100110";
		Trees_din <= x"00046410";
		wait for Clk_period;
		Addr <=  "00001011100111";
		Trees_din <= x"18004608";
		wait for Clk_period;
		Addr <=  "00001011101000";
		Trees_din <= x"1900a004";
		wait for Clk_period;
		Addr <=  "00001011101001";
		Trees_din <= x"ffd70bc5";
		wait for Clk_period;
		Addr <=  "00001011101010";
		Trees_din <= x"00230bc5";
		wait for Clk_period;
		Addr <=  "00001011101011";
		Trees_din <= x"1e007804";
		wait for Clk_period;
		Addr <=  "00001011101100";
		Trees_din <= x"00620bc5";
		wait for Clk_period;
		Addr <=  "00001011101101";
		Trees_din <= x"000a0bc5";
		wait for Clk_period;
		Addr <=  "00001011101110";
		Trees_din <= x"06023204";
		wait for Clk_period;
		Addr <=  "00001011101111";
		Trees_din <= x"ffaa0bc5";
		wait for Clk_period;
		Addr <=  "00001011110000";
		Trees_din <= x"00070bc5";
		wait for Clk_period;
		Addr <=  "00001011110001";
		Trees_din <= x"06f9ca04";
		wait for Clk_period;
		Addr <=  "00001011110010";
		Trees_din <= x"ff890bf9";
		wait for Clk_period;
		Addr <=  "00001011110011";
		Trees_din <= x"06091b10";
		wait for Clk_period;
		Addr <=  "00001011110100";
		Trees_din <= x"0d003004";
		wait for Clk_period;
		Addr <=  "00001011110101";
		Trees_din <= x"00300bf9";
		wait for Clk_period;
		Addr <=  "00001011110110";
		Trees_din <= x"14014604";
		wait for Clk_period;
		Addr <=  "00001011110111";
		Trees_din <= x"ffa50bf9";
		wait for Clk_period;
		Addr <=  "00001011111000";
		Trees_din <= x"16022d04";
		wait for Clk_period;
		Addr <=  "00001011111001";
		Trees_din <= x"ffd60bf9";
		wait for Clk_period;
		Addr <=  "00001011111010";
		Trees_din <= x"00220bf9";
		wait for Clk_period;
		Addr <=  "00001011111011";
		Trees_din <= x"0e01d204";
		wait for Clk_period;
		Addr <=  "00001011111100";
		Trees_din <= x"00530bf9";
		wait for Clk_period;
		Addr <=  "00001011111101";
		Trees_din <= x"000c0bf9";
		wait for Clk_period;
		Addr <=  "00001011111110";
		Trees_din <= x"06f9ca04";
		wait for Clk_period;
		Addr <=  "00001011111111";
		Trees_din <= x"ff8c0c25";
		wait for Clk_period;
		Addr <=  "00001100000000";
		Trees_din <= x"01070110";
		wait for Clk_period;
		Addr <=  "00001100000001";
		Trees_din <= x"06091b0c";
		wait for Clk_period;
		Addr <=  "00001100000010";
		Trees_din <= x"13f96104";
		wait for Clk_period;
		Addr <=  "00001100000011";
		Trees_din <= x"00310c25";
		wait for Clk_period;
		Addr <=  "00001100000100";
		Trees_din <= x"0e024004";
		wait for Clk_period;
		Addr <=  "00001100000101";
		Trees_din <= x"ffbc0c25";
		wait for Clk_period;
		Addr <=  "00001100000110";
		Trees_din <= x"001a0c25";
		wait for Clk_period;
		Addr <=  "00001100000111";
		Trees_din <= x"00520c25";
		wait for Clk_period;
		Addr <=  "00001100001000";
		Trees_din <= x"ffc00c25";
		wait for Clk_period;
		Addr <=  "00001100001001";
		Trees_din <= x"06f9ca04";
		wait for Clk_period;
		Addr <=  "00001100001010";
		Trees_din <= x"ff900c59";
		wait for Clk_period;
		Addr <=  "00001100001011";
		Trees_din <= x"00046410";
		wait for Clk_period;
		Addr <=  "00001100001100";
		Trees_din <= x"18004408";
		wait for Clk_period;
		Addr <=  "00001100001101";
		Trees_din <= x"03013f04";
		wait for Clk_period;
		Addr <=  "00001100001110";
		Trees_din <= x"00280c59";
		wait for Clk_period;
		Addr <=  "00001100001111";
		Trees_din <= x"ffd50c59";
		wait for Clk_period;
		Addr <=  "00001100010000";
		Trees_din <= x"1a00b404";
		wait for Clk_period;
		Addr <=  "00001100010001";
		Trees_din <= x"00020c59";
		wait for Clk_period;
		Addr <=  "00001100010010";
		Trees_din <= x"005c0c59";
		wait for Clk_period;
		Addr <=  "00001100010011";
		Trees_din <= x"02ffb904";
		wait for Clk_period;
		Addr <=  "00001100010100";
		Trees_din <= x"00030c59";
		wait for Clk_period;
		Addr <=  "00001100010101";
		Trees_din <= x"ffb10c59";
		wait for Clk_period;
		Addr <=  "00001100010110";
		Trees_din <= x"06ffc308";
		wait for Clk_period;
		Addr <=  "00001100010111";
		Trees_din <= x"02fe2704";
		wait for Clk_period;
		Addr <=  "00001100011000";
		Trees_din <= x"000a0c85";
		wait for Clk_period;
		Addr <=  "00001100011001";
		Trees_din <= x"ff8c0c85";
		wait for Clk_period;
		Addr <=  "00001100011010";
		Trees_din <= x"06091b0c";
		wait for Clk_period;
		Addr <=  "00001100011011";
		Trees_din <= x"0c028d08";
		wait for Clk_period;
		Addr <=  "00001100011100";
		Trees_din <= x"0b027504";
		wait for Clk_period;
		Addr <=  "00001100011101";
		Trees_din <= x"ffff0c85";
		wait for Clk_period;
		Addr <=  "00001100011110";
		Trees_din <= x"ffbd0c85";
		wait for Clk_period;
		Addr <=  "00001100011111";
		Trees_din <= x"00290c85";
		wait for Clk_period;
		Addr <=  "00001100100000";
		Trees_din <= x"003b0c85";
		wait for Clk_period;
		Addr <=  "00001100100001";
		Trees_din <= x"06f9ca04";
		wait for Clk_period;
		Addr <=  "00001100100010";
		Trees_din <= x"ff980cb1";
		wait for Clk_period;
		Addr <=  "00001100100011";
		Trees_din <= x"13f96908";
		wait for Clk_period;
		Addr <=  "00001100100100";
		Trees_din <= x"02fe0104";
		wait for Clk_period;
		Addr <=  "00001100100101";
		Trees_din <= x"004b0cb1";
		wait for Clk_period;
		Addr <=  "00001100100110";
		Trees_din <= x"00050cb1";
		wait for Clk_period;
		Addr <=  "00001100100111";
		Trees_din <= x"16007904";
		wait for Clk_period;
		Addr <=  "00001100101000";
		Trees_din <= x"00200cb1";
		wait for Clk_period;
		Addr <=  "00001100101001";
		Trees_din <= x"09005704";
		wait for Clk_period;
		Addr <=  "00001100101010";
		Trees_din <= x"ffbc0cb1";
		wait for Clk_period;
		Addr <=  "00001100101011";
		Trees_din <= x"00080cb1";
		wait for Clk_period;
		Addr <=  "00001100101100";
		Trees_din <= x"06ffc308";
		wait for Clk_period;
		Addr <=  "00001100101101";
		Trees_din <= x"12fec504";
		wait for Clk_period;
		Addr <=  "00001100101110";
		Trees_din <= x"00050cdd";
		wait for Clk_period;
		Addr <=  "00001100101111";
		Trees_din <= x"ff940cdd";
		wait for Clk_period;
		Addr <=  "00001100110000";
		Trees_din <= x"06091b0c";
		wait for Clk_period;
		Addr <=  "00001100110001";
		Trees_din <= x"03fbbc04";
		wait for Clk_period;
		Addr <=  "00001100110010";
		Trees_din <= x"002b0cdd";
		wait for Clk_period;
		Addr <=  "00001100110011";
		Trees_din <= x"0c015d04";
		wait for Clk_period;
		Addr <=  "00001100110100";
		Trees_din <= x"fffe0cdd";
		wait for Clk_period;
		Addr <=  "00001100110101";
		Trees_din <= x"ffc00cdd";
		wait for Clk_period;
		Addr <=  "00001100110110";
		Trees_din <= x"00380cdd";
		wait for Clk_period;
		Addr <=  "00001100110111";
		Trees_din <= x"06ffc308";
		wait for Clk_period;
		Addr <=  "00001100111000";
		Trees_din <= x"12fec504";
		wait for Clk_period;
		Addr <=  "00001100111001";
		Trees_din <= x"00030d09";
		wait for Clk_period;
		Addr <=  "00001100111010";
		Trees_din <= x"ff980d09";
		wait for Clk_period;
		Addr <=  "00001100111011";
		Trees_din <= x"04f47104";
		wait for Clk_period;
		Addr <=  "00001100111100";
		Trees_din <= x"ffdd0d09";
		wait for Clk_period;
		Addr <=  "00001100111101";
		Trees_din <= x"03fbbc04";
		wait for Clk_period;
		Addr <=  "00001100111110";
		Trees_din <= x"00410d09";
		wait for Clk_period;
		Addr <=  "00001100111111";
		Trees_din <= x"05fb9304";
		wait for Clk_period;
		Addr <=  "00001101000000";
		Trees_din <= x"00220d09";
		wait for Clk_period;
		Addr <=  "00001101000001";
		Trees_din <= x"ffd80d09";
		wait for Clk_period;
		Addr <=  "00001101000010";
		Trees_din <= x"06f9ca04";
		wait for Clk_period;
		Addr <=  "00001101000011";
		Trees_din <= x"ffa30d2d";
		wait for Clk_period;
		Addr <=  "00001101000100";
		Trees_din <= x"02002408";
		wait for Clk_period;
		Addr <=  "00001101000101";
		Trees_din <= x"0d017a04";
		wait for Clk_period;
		Addr <=  "00001101000110";
		Trees_din <= x"003e0d2d";
		wait for Clk_period;
		Addr <=  "00001101000111";
		Trees_din <= x"fff20d2d";
		wait for Clk_period;
		Addr <=  "00001101001000";
		Trees_din <= x"16024704";
		wait for Clk_period;
		Addr <=  "00001101001001";
		Trees_din <= x"ffff0d2d";
		wait for Clk_period;
		Addr <=  "00001101001010";
		Trees_din <= x"ffcb0d2d";
		wait for Clk_period;
		Addr <=  "00001101001011";
		Trees_din <= x"06091b10";
		wait for Clk_period;
		Addr <=  "00001101001100";
		Trees_din <= x"13f96104";
		wait for Clk_period;
		Addr <=  "00001101001101";
		Trees_din <= x"000c0d51";
		wait for Clk_period;
		Addr <=  "00001101001110";
		Trees_din <= x"0600ad04";
		wait for Clk_period;
		Addr <=  "00001101001111";
		Trees_din <= x"ff9b0d51";
		wait for Clk_period;
		Addr <=  "00001101010000";
		Trees_din <= x"1401e904";
		wait for Clk_period;
		Addr <=  "00001101010001";
		Trees_din <= x"ffcf0d51";
		wait for Clk_period;
		Addr <=  "00001101010010";
		Trees_din <= x"001a0d51";
		wait for Clk_period;
		Addr <=  "00001101010011";
		Trees_din <= x"00350d51";
		wait for Clk_period;
		Addr <=  "00001101010100";
		Trees_din <= x"06091b0c";
		wait for Clk_period;
		Addr <=  "00001101010101";
		Trees_din <= x"0003aa08";
		wait for Clk_period;
		Addr <=  "00001101010110";
		Trees_din <= x"1004b404";
		wait for Clk_period;
		Addr <=  "00001101010111";
		Trees_din <= x"ffda0d6d";
		wait for Clk_period;
		Addr <=  "00001101011000";
		Trees_din <= x"001d0d6d";
		wait for Clk_period;
		Addr <=  "00001101011001";
		Trees_din <= x"ffb00d6d";
		wait for Clk_period;
		Addr <=  "00001101011010";
		Trees_din <= x"00320d6d";
		wait for Clk_period;
		Addr <=  "00001101011011";
		Trees_din <= x"06f9ca04";
		wait for Clk_period;
		Addr <=  "00001101011100";
		Trees_din <= x"ffad0d91";
		wait for Clk_period;
		Addr <=  "00001101011101";
		Trees_din <= x"01060b0c";
		wait for Clk_period;
		Addr <=  "00001101011110";
		Trees_din <= x"1d004808";
		wait for Clk_period;
		Addr <=  "00001101011111";
		Trees_din <= x"18004204";
		wait for Clk_period;
		Addr <=  "00001101100000";
		Trees_din <= x"ffff0d91";
		wait for Clk_period;
		Addr <=  "00001101100001";
		Trees_din <= x"00420d91";
		wait for Clk_period;
		Addr <=  "00001101100010";
		Trees_din <= x"fff50d91";
		wait for Clk_period;
		Addr <=  "00001101100011";
		Trees_din <= x"ffd20d91";
		wait for Clk_period;
		Addr <=  "00001101100100";
		Trees_din <= x"06091b10";
		wait for Clk_period;
		Addr <=  "00001101100101";
		Trees_din <= x"0d003004";
		wait for Clk_period;
		Addr <=  "00001101100110";
		Trees_din <= x"00150db5";
		wait for Clk_period;
		Addr <=  "00001101100111";
		Trees_din <= x"06fee904";
		wait for Clk_period;
		Addr <=  "00001101101000";
		Trees_din <= x"ffa60db5";
		wait for Clk_period;
		Addr <=  "00001101101001";
		Trees_din <= x"0c02a404";
		wait for Clk_period;
		Addr <=  "00001101101010";
		Trees_din <= x"ffd60db5";
		wait for Clk_period;
		Addr <=  "00001101101011";
		Trees_din <= x"00170db5";
		wait for Clk_period;
		Addr <=  "00001101101100";
		Trees_din <= x"00300db5";
		wait for Clk_period;
		Addr <=  "00001101101101";
		Trees_din <= x"0003e50c";
		wait for Clk_period;
		Addr <=  "00001101101110";
		Trees_din <= x"18004404";
		wait for Clk_period;
		Addr <=  "00001101101111";
		Trees_din <= x"fff20dd9";
		wait for Clk_period;
		Addr <=  "00001101110000";
		Trees_din <= x"1a00b404";
		wait for Clk_period;
		Addr <=  "00001101110001";
		Trees_din <= x"fffb0dd9";
		wait for Clk_period;
		Addr <=  "00001101110010";
		Trees_din <= x"00440dd9";
		wait for Clk_period;
		Addr <=  "00001101110011";
		Trees_din <= x"02004a04";
		wait for Clk_period;
		Addr <=  "00001101110100";
		Trees_din <= x"fff70dd9";
		wait for Clk_period;
		Addr <=  "00001101110101";
		Trees_din <= x"ffb00dd9";
		wait for Clk_period;
		Addr <=  "00001101110110";
		Trees_din <= x"06ffc304";
		wait for Clk_period;
		Addr <=  "00001101110111";
		Trees_din <= x"ffc60df5";
		wait for Clk_period;
		Addr <=  "00001101111000";
		Trees_din <= x"1900a008";
		wait for Clk_period;
		Addr <=  "00001101111001";
		Trees_din <= x"11028704";
		wait for Clk_period;
		Addr <=  "00001101111010";
		Trees_din <= x"ffd90df5";
		wait for Clk_period;
		Addr <=  "00001101111011";
		Trees_din <= x"00220df5";
		wait for Clk_period;
		Addr <=  "00001101111100";
		Trees_din <= x"00340df5";
		wait for Clk_period;
		Addr <=  "00001101111101";
		Trees_din <= x"0004640c";
		wait for Clk_period;
		Addr <=  "00001101111110";
		Trees_din <= x"18004404";
		wait for Clk_period;
		Addr <=  "00001101111111";
		Trees_din <= x"fff30e11";
		wait for Clk_period;
		Addr <=  "00001110000000";
		Trees_din <= x"1a00b404";
		wait for Clk_period;
		Addr <=  "00001110000001";
		Trees_din <= x"00010e11";
		wait for Clk_period;
		Addr <=  "00001110000010";
		Trees_din <= x"00410e11";
		wait for Clk_period;
		Addr <=  "00001110000011";
		Trees_din <= x"ffca0e11";
		wait for Clk_period;
		Addr <=  "00001110000100";
		Trees_din <= x"06091b0c";
		wait for Clk_period;
		Addr <=  "00001110000101";
		Trees_din <= x"13f96104";
		wait for Clk_period;
		Addr <=  "00001110000110";
		Trees_din <= x"00120e2d";
		wait for Clk_period;
		Addr <=  "00001110000111";
		Trees_din <= x"06054004";
		wait for Clk_period;
		Addr <=  "00001110001000";
		Trees_din <= x"ffb50e2d";
		wait for Clk_period;
		Addr <=  "00001110001001";
		Trees_din <= x"00040e2d";
		wait for Clk_period;
		Addr <=  "00001110001010";
		Trees_din <= x"00300e2d";
		wait for Clk_period;
		Addr <=  "00001110001011";
		Trees_din <= x"0107010c";
		wait for Clk_period;
		Addr <=  "00001110001100";
		Trees_din <= x"05f9ce04";
		wait for Clk_period;
		Addr <=  "00001110001101";
		Trees_din <= x"002f0e49";
		wait for Clk_period;
		Addr <=  "00001110001110";
		Trees_din <= x"08008504";
		wait for Clk_period;
		Addr <=  "00001110001111";
		Trees_din <= x"00190e49";
		wait for Clk_period;
		Addr <=  "00001110010000";
		Trees_din <= x"ffda0e49";
		wait for Clk_period;
		Addr <=  "00001110010001";
		Trees_din <= x"ffc00e49";
		wait for Clk_period;
		Addr <=  "00001110010010";
		Trees_din <= x"02002408";
		wait for Clk_period;
		Addr <=  "00001110010011";
		Trees_din <= x"0d017504";
		wait for Clk_period;
		Addr <=  "00001110010100";
		Trees_din <= x"002e0e65";
		wait for Clk_period;
		Addr <=  "00001110010101";
		Trees_din <= x"fff30e65";
		wait for Clk_period;
		Addr <=  "00001110010110";
		Trees_din <= x"16024704";
		wait for Clk_period;
		Addr <=  "00001110010111";
		Trees_din <= x"fff50e65";
		wait for Clk_period;
		Addr <=  "00001110011000";
		Trees_din <= x"ffc90e65";
		wait for Clk_period;
		Addr <=  "00001110011001";
		Trees_din <= x"06054008";
		wait for Clk_period;
		Addr <=  "00001110011010";
		Trees_din <= x"13f96104";
		wait for Clk_period;
		Addr <=  "00001110011011";
		Trees_din <= x"00140e81";
		wait for Clk_period;
		Addr <=  "00001110011100";
		Trees_din <= x"ffb90e81";
		wait for Clk_period;
		Addr <=  "00001110011101";
		Trees_din <= x"0c01cb04";
		wait for Clk_period;
		Addr <=  "00001110011110";
		Trees_din <= x"00330e81";
		wait for Clk_period;
		Addr <=  "00001110011111";
		Trees_din <= x"fffa0e81";
		wait for Clk_period;
		Addr <=  "00001110100000";
		Trees_din <= x"06091b0c";
		wait for Clk_period;
		Addr <=  "00001110100001";
		Trees_din <= x"0d003004";
		wait for Clk_period;
		Addr <=  "00001110100010";
		Trees_din <= x"00140e9d";
		wait for Clk_period;
		Addr <=  "00001110100011";
		Trees_din <= x"0f00ff04";
		wait for Clk_period;
		Addr <=  "00001110100100";
		Trees_din <= x"ffb70e9d";
		wait for Clk_period;
		Addr <=  "00001110100101";
		Trees_din <= x"fff90e9d";
		wait for Clk_period;
		Addr <=  "00001110100110";
		Trees_din <= x"002c0e9d";
		wait for Clk_period;
		Addr <=  "00001110100111";
		Trees_din <= x"00046408";
		wait for Clk_period;
		Addr <=  "00001110101000";
		Trees_din <= x"18004404";
		wait for Clk_period;
		Addr <=  "00001110101001";
		Trees_din <= x"fff40eb1";
		wait for Clk_period;
		Addr <=  "00001110101010";
		Trees_din <= x"00280eb1";
		wait for Clk_period;
		Addr <=  "00001110101011";
		Trees_din <= x"ffd20eb1";
		wait for Clk_period;
		Addr <=  "00001110101100";
		Trees_din <= x"06091b0c";
		wait for Clk_period;
		Addr <=  "00001110101101";
		Trees_din <= x"0d003004";
		wait for Clk_period;
		Addr <=  "00001110101110";
		Trees_din <= x"00120ecd";
		wait for Clk_period;
		Addr <=  "00001110101111";
		Trees_din <= x"0f00ff04";
		wait for Clk_period;
		Addr <=  "00001110110000";
		Trees_din <= x"ffbb0ecd";
		wait for Clk_period;
		Addr <=  "00001110110001";
		Trees_din <= x"fffa0ecd";
		wait for Clk_period;
		Addr <=  "00001110110010";
		Trees_din <= x"00290ecd";
		wait for Clk_period;
		Addr <=  "00001110110011";
		Trees_din <= x"02002408";
		wait for Clk_period;
		Addr <=  "00001110110100";
		Trees_din <= x"0d019304";
		wait for Clk_period;
		Addr <=  "00001110110101";
		Trees_din <= x"00280ee1";
		wait for Clk_period;
		Addr <=  "00001110110110";
		Trees_din <= x"fff50ee1";
		wait for Clk_period;
		Addr <=  "00001110110111";
		Trees_din <= x"ffd90ee1";
		wait for Clk_period;
		Addr <=  "00001110111000";
		Trees_din <= x"00046408";
		wait for Clk_period;
		Addr <=  "00001110111001";
		Trees_din <= x"18004404";
		wait for Clk_period;
		Addr <=  "00001110111010";
		Trees_din <= x"fff60ef5";
		wait for Clk_period;
		Addr <=  "00001110111011";
		Trees_din <= x"00250ef5";
		wait for Clk_period;
		Addr <=  "00001110111100";
		Trees_din <= x"ffd60ef5";
		wait for Clk_period;
		Addr <=  "00001110111101";
		Trees_din <= x"06ffc304";
		wait for Clk_period;
		Addr <=  "00001110111110";
		Trees_din <= x"ffd40f11";
		wait for Clk_period;
		Addr <=  "00001110111111";
		Trees_din <= x"1900a008";
		wait for Clk_period;
		Addr <=  "00001111000000";
		Trees_din <= x"11028404";
		wait for Clk_period;
		Addr <=  "00001111000001";
		Trees_din <= x"ffe10f11";
		wait for Clk_period;
		Addr <=  "00001111000010";
		Trees_din <= x"00140f11";
		wait for Clk_period;
		Addr <=  "00001111000011";
		Trees_din <= x"00330f11";
		wait for Clk_period;
		Addr <=  "00001111000100";
		Trees_din <= x"13f96904";
		wait for Clk_period;
		Addr <=  "00001111000101";
		Trees_din <= x"00210f25";
		wait for Clk_period;
		Addr <=  "00001111000110";
		Trees_din <= x"06054004";
		wait for Clk_period;
		Addr <=  "00001111000111";
		Trees_din <= x"ffc70f25";
		wait for Clk_period;
		Addr <=  "00001111001000";
		Trees_din <= x"000e0f25";
		wait for Clk_period;
		Addr <=  "00001111001001";
		Trees_din <= x"0000001f";
		wait for Clk_period;

        -- Reset valid flag
        Valid_node <= '0';
        wait for Clk_period; 
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001000100011100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010011001100";
        wait for Clk_period; 
        Features_din <= "0000011010100101";
        wait for Clk_period; 
        Features_din <= "1111100111011011";
        wait for Clk_period; 
        Features_din <= "1111110000001010";
        wait for Clk_period; 
        Features_din <= "0000001010001101";
        wait for Clk_period; 
        Features_din <= "1111010001011001";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000100111011";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "1111101100000001";
        wait for Clk_period; 
        Features_din <= "1111100101001101";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001000101101";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000010100011100";
        wait for Clk_period; 
        Features_din <= "0000001010100110";
        wait for Clk_period; 
        Features_din <= "0000001000001101";
        wait for Clk_period; 
        Features_din <= "1111111110110110";
        wait for Clk_period; 
        Features_din <= "0000000011011110";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000001100010101";
        wait for Clk_period; 
        Features_din <= "0000000100010010";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000110111110111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001010001001000";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "1111000100111111";
        wait for Clk_period; 
        Features_din <= "1111100101101010";
        wait for Clk_period; 
        Features_din <= "1111111010101111";
        wait for Clk_period; 
        Features_din <= "1111000110100011";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000001010001000";
        wait for Clk_period; 
        Features_din <= "0000001010001000";
        wait for Clk_period; 
        Features_din <= "0000000110001110";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111100110100101";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000001010001000";
        wait for Clk_period; 
        Features_din <= "0000001010001000";
        wait for Clk_period; 
        Features_din <= "0000001010001000";
        wait for Clk_period; 
        Features_din <= "1111100110110101";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000000011111100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001011010001101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000100111100111";
        wait for Clk_period; 
        Features_din <= "1111101110010111";
        wait for Clk_period; 
        Features_din <= "1111010111111110";
        wait for Clk_period; 
        Features_din <= "1111110000001111";
        wait for Clk_period; 
        Features_din <= "1111110001001111";
        wait for Clk_period; 
        Features_din <= "1111000110100101";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000000011110010";
        wait for Clk_period; 
        Features_din <= "0000001000100111";
        wait for Clk_period; 
        Features_din <= "0000000100100101";
        wait for Clk_period; 
        Features_din <= "0000010100100111";
        wait for Clk_period; 
        Features_din <= "0000000011101101";
        wait for Clk_period; 
        Features_din <= "1111100010000111";
        wait for Clk_period; 
        Features_din <= "0000000110101011";
        wait for Clk_period; 
        Features_din <= "1111111001010111";
        wait for Clk_period; 
        Features_din <= "1111110101011001";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000000110110011";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "0000000011101001";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010010111110010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001011010001";
        wait for Clk_period; 
        Features_din <= "1110110101000111";
        wait for Clk_period; 
        Features_din <= "1110111101001011";
        wait for Clk_period; 
        Features_din <= "1111101100100000";
        wait for Clk_period; 
        Features_din <= "1111011110111101";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000111111100";
        wait for Clk_period; 
        Features_din <= "0000010100110001";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "0000001010111010";
        wait for Clk_period; 
        Features_din <= "1111111001000011";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000010010100111";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "1111111000000011";
        wait for Clk_period; 
        Features_din <= "1111100011010000";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001011010011";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111101101001110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111000111001";
        wait for Clk_period; 
        Features_din <= "0000101001111100";
        wait for Clk_period; 
        Features_din <= "1111111011001011";
        wait for Clk_period; 
        Features_din <= "1111111110010011";
        wait for Clk_period; 
        Features_din <= "0000100000001010";
        wait for Clk_period; 
        Features_din <= "1111001011100001";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000000100001000";
        wait for Clk_period; 
        Features_din <= "0000000101011100";
        wait for Clk_period; 
        Features_din <= "1111011011111011";
        wait for Clk_period; 
        Features_din <= "0000000110001010";
        wait for Clk_period; 
        Features_din <= "0000000100011001";
        wait for Clk_period; 
        Features_din <= "1111111010011101";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000110110011";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001011000010001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111101001001000";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "1111100010000010";
        wait for Clk_period; 
        Features_din <= "1111110111000000";
        wait for Clk_period; 
        Features_din <= "1111111100101000";
        wait for Clk_period; 
        Features_din <= "1111111010101100";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000000111001000";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111111001001010";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010100000000";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "1111110111110101";
        wait for Clk_period; 
        Features_din <= "1111100010100000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "0000000011000000";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000010001010101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010100101010";
        wait for Clk_period; 
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "1111100000001100";
        wait for Clk_period; 
        Features_din <= "1111011000101000";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000100001010";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000100110001";
        wait for Clk_period; 
        Features_din <= "0000010101001001";
        wait for Clk_period; 
        Features_din <= "0000001100010001";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "1111110100011110";
        wait for Clk_period; 
        Features_din <= "0000001000110010";
        wait for Clk_period; 
        Features_din <= "0000010100100011";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "1111111001100110";
        wait for Clk_period; 
        Features_din <= "1111100101000110";
        wait for Clk_period; 
        Features_din <= "0000000111011111";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "0000000101010110";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "0000000011100101";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001000010110111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111110010110100";
        wait for Clk_period; 
        Features_din <= "0000000110011001";
        wait for Clk_period; 
        Features_din <= "1111100100011010";
        wait for Clk_period; 
        Features_din <= "1111101001000111";
        wait for Clk_period; 
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "1111110011100111";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000111011011";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111101010110001";
        wait for Clk_period; 
        Features_din <= "1111110010000011";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000000100101000";
        wait for Clk_period; 
        Features_din <= "0000011001000111";
        wait for Clk_period; 
        Features_din <= "0000001000011100";
        wait for Clk_period; 
        Features_din <= "0000010010000110";
        wait for Clk_period; 
        Features_din <= "0000000101000011";
        wait for Clk_period; 
        Features_din <= "1111111111101100";
        wait for Clk_period; 
        Features_din <= "1111110011001111";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000000010111111";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010100111001011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "1111101111011110";
        wait for Clk_period; 
        Features_din <= "1110101100001000";
        wait for Clk_period; 
        Features_din <= "1111000011011010";
        wait for Clk_period; 
        Features_din <= "1111101111100011";
        wait for Clk_period; 
        Features_din <= "1111010100000100";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000101111100";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000000011001000";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111100111110011";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "1111100101101001";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000011011101";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001011101101001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000100011101110";
        wait for Clk_period; 
        Features_din <= "0000110000011000";
        wait for Clk_period; 
        Features_din <= "1111000011010000";
        wait for Clk_period; 
        Features_din <= "1111101101111100";
        wait for Clk_period; 
        Features_din <= "1111011101111001";
        wait for Clk_period; 
        Features_din <= "1111010110010110";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000001001110100";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111100000010001";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001000100010";
        wait for Clk_period; 
        Features_din <= "0000000101111111";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000010011111010";
        wait for Clk_period; 
        Features_din <= "0000000111010100";
        wait for Clk_period; 
        Features_din <= "1111111110101100";
        wait for Clk_period; 
        Features_din <= "1111110101000100";
        wait for Clk_period; 
        Features_din <= "0000000101111100";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000011001011";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000111001011101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000000011110010";
        wait for Clk_period; 
        Features_din <= "0000001000000110";
        wait for Clk_period; 
        Features_din <= "1111110010011111";
        wait for Clk_period; 
        Features_din <= "1111101100100100";
        wait for Clk_period; 
        Features_din <= "1111111000010001";
        wait for Clk_period; 
        Features_din <= "1111010010110110";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000011001001";
        wait for Clk_period; 
        Features_din <= "1111111000000111";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "1111111110000001";
        wait for Clk_period; 
        Features_din <= "1111100000001110";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001111011001011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011010010101";
        wait for Clk_period; 
        Features_din <= "1111111100111011";
        wait for Clk_period; 
        Features_din <= "1111000101101110";
        wait for Clk_period; 
        Features_din <= "1111001101010010";
        wait for Clk_period; 
        Features_din <= "1111110011011001";
        wait for Clk_period; 
        Features_din <= "1111101011111101";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000101000100";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111111101000110";
        wait for Clk_period; 
        Features_din <= "1111101101100010";
        wait for Clk_period; 
        Features_din <= "0000001001011001";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "1111101000001000";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000000100111110";
        wait for Clk_period; 
        Features_din <= "0000011000100001";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "0000000011001000";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010111110010101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111011111000011";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "1111011101001110";
        wait for Clk_period; 
        Features_din <= "1111010001100011";
        wait for Clk_period; 
        Features_din <= "1111101001000110";
        wait for Clk_period; 
        Features_din <= "1111011110001001";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000001010010000";
        wait for Clk_period; 
        Features_din <= "0000010010110000";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "0000001100101001";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "1111011101000001";
        wait for Clk_period; 
        Features_din <= "0000000101111000";
        wait for Clk_period; 
        Features_din <= "0000000100101000";
        wait for Clk_period; 
        Features_din <= "1111111000111110";
        wait for Clk_period; 
        Features_din <= "0000001001110000";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000101110110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001001011100";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000011000001010";
        wait for Clk_period; 
        Features_din <= "0000000110010100";
        wait for Clk_period; 
        Features_din <= "1111110011111110";
        wait for Clk_period; 
        Features_din <= "1111110100001001";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000011111000";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111101100001100";
        wait for Clk_period; 
        Features_din <= "0000010101011111";
        wait for Clk_period; 
        Features_din <= "0000000110111000";
        wait for Clk_period; 
        Features_din <= "0000001010010010";
        wait for Clk_period; 
        Features_din <= "0000000111010111";
        wait for Clk_period; 
        Features_din <= "0000000100001001";
        wait for Clk_period; 
        Features_din <= "1111100101011000";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "0000001000100100";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "0000000100000111";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001010111000";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010011100101100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010101011010";
        wait for Clk_period; 
        Features_din <= "1111110101011110";
        wait for Clk_period; 
        Features_din <= "1110101111100101";
        wait for Clk_period; 
        Features_din <= "1111010111100111";
        wait for Clk_period; 
        Features_din <= "1111010010101110";
        wait for Clk_period; 
        Features_din <= "1111011101100000";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000010101100";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111110011001111";
        wait for Clk_period; 
        Features_din <= "1111101100010110";
        wait for Clk_period; 
        Features_din <= "0000000111001001";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000000011001000";
        wait for Clk_period; 
        Features_din <= "1111101010110100";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000000110001001";
        wait for Clk_period; 
        Features_din <= "0000000100111000";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001000110001001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000100001000010";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "1111101011001101";
        wait for Clk_period; 
        Features_din <= "1111011001011000";
        wait for Clk_period; 
        Features_din <= "1111010100100001";
        wait for Clk_period; 
        Features_din <= "1111111000111110";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000110010110";
        wait for Clk_period; 
        Features_din <= "0000010100100100";
        wait for Clk_period; 
        Features_din <= "0000000100011100";
        wait for Clk_period; 
        Features_din <= "0000001010110000";
        wait for Clk_period; 
        Features_din <= "1111110110100110";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000010100100100";
        wait for Clk_period; 
        Features_din <= "1111111010101000";
        wait for Clk_period; 
        Features_din <= "1111111010111011";
        wait for Clk_period; 
        Features_din <= "1111100100011000";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001011110100";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0011001001001001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000110111000000";
        wait for Clk_period; 
        Features_din <= "1111010101101111";
        wait for Clk_period; 
        Features_din <= "1111000000011011";
        wait for Clk_period; 
        Features_din <= "1110111101111011";
        wait for Clk_period; 
        Features_din <= "1111001100001001";
        wait for Clk_period; 
        Features_din <= "1111000011010111";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000000111011000";
        wait for Clk_period; 
        Features_din <= "0000000110010111";
        wait for Clk_period; 
        Features_din <= "1111100110000011";
        wait for Clk_period; 
        Features_din <= "0000001011101101";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "1111100111010111";
        wait for Clk_period; 
        Features_din <= "0000001011000011";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "0000001000000011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010101110111100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000110010011100";
        wait for Clk_period; 
        Features_din <= "0000001011101101";
        wait for Clk_period; 
        Features_din <= "1110110010010001";
        wait for Clk_period; 
        Features_din <= "1111011101011000";
        wait for Clk_period; 
        Features_din <= "1111110100000101";
        wait for Clk_period; 
        Features_din <= "1111011010011011";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000111010000";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111101101111110";
        wait for Clk_period; 
        Features_din <= "0000011100010001";
        wait for Clk_period; 
        Features_din <= "0000001001000101";
        wait for Clk_period; 
        Features_din <= "0000001010100110";
        wait for Clk_period; 
        Features_din <= "1111111101100111";
        wait for Clk_period; 
        Features_din <= "0000000101001110";
        wait for Clk_period; 
        Features_din <= "1111110110100000";
        wait for Clk_period; 
        Features_din <= "1111101101101101";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000000101100100";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000001100000110";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000111101000000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "1111101110001110";
        wait for Clk_period; 
        Features_din <= "1111101101111100";
        wait for Clk_period; 
        Features_din <= "1111110001111100";
        wait for Clk_period; 
        Features_din <= "1111101110100100";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000000011110011";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "1111110110101011";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "1111011111101110";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001000000100";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000011000100";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110110010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000100000001010";
        wait for Clk_period; 
        Features_din <= "1111111110010000";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "0000100111111011";
        wait for Clk_period; 
        Features_din <= "1111011101010010";
        wait for Clk_period; 
        Features_din <= "1111001110101110";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000101111110";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "1111100111111000";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001011111010";
        wait for Clk_period; 
        Features_din <= "0000001000110101";
        wait for Clk_period; 
        Features_din <= "0000000100010111";
        wait for Clk_period; 
        Features_din <= "1111100111011000";
        wait for Clk_period; 
        Features_din <= "0000001001011100";
        wait for Clk_period; 
        Features_din <= "0000001100001101";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000001000101100";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000100111101";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000010101101";
        wait for Clk_period; 
        Features_din <= "0000000011100000";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001100111001110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010011000100";
        wait for Clk_period; 
        Features_din <= "1111110010101001";
        wait for Clk_period; 
        Features_din <= "1111011011101001";
        wait for Clk_period; 
        Features_din <= "1111111010000111";
        wait for Clk_period; 
        Features_din <= "1111111000000000";
        wait for Clk_period; 
        Features_din <= "1111100101101000";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111101100101111";
        wait for Clk_period; 
        Features_din <= "1111100111011110";
        wait for Clk_period; 
        Features_din <= "0000001100001100";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000000111001111";
        wait for Clk_period; 
        Features_din <= "0000000100111011";
        wait for Clk_period; 
        Features_din <= "0000011001101011";
        wait for Clk_period; 
        Features_din <= "0000001000101010";
        wait for Clk_period; 
        Features_din <= "0000000101000010";
        wait for Clk_period; 
        Features_din <= "1111111101001101";
        wait for Clk_period; 
        Features_din <= "0000001000111000";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000001001001000";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000000010111111";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001000011011000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001010010000";
        wait for Clk_period; 
        Features_din <= "0001000011000101";
        wait for Clk_period; 
        Features_din <= "1111011110001100";
        wait for Clk_period; 
        Features_din <= "1111010110001010";
        wait for Clk_period; 
        Features_din <= "1111101011111000";
        wait for Clk_period; 
        Features_din <= "1111000111101001";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000011000101111";
        wait for Clk_period; 
        Features_din <= "1111111011110010";
        wait for Clk_period; 
        Features_din <= "0000001000111100";
        wait for Clk_period; 
        Features_din <= "0000000101011011";
        wait for Clk_period; 
        Features_din <= "1111110110001011";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000011000000001";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "1111110011111011";
        wait for Clk_period; 
        Features_din <= "1111101110000101";
        wait for Clk_period; 
        Features_din <= "0000000111100101";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "0000001001000011";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001111101111000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010111110011";
        wait for Clk_period; 
        Features_din <= "1111111110010001";
        wait for Clk_period; 
        Features_din <= "1111001010110010";
        wait for Clk_period; 
        Features_din <= "1111010000110100";
        wait for Clk_period; 
        Features_din <= "1111101011111000";
        wait for Clk_period; 
        Features_din <= "1111100001000010";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111011111011100";
        wait for Clk_period; 
        Features_din <= "0000010011111100";
        wait for Clk_period; 
        Features_din <= "0000001010101111";
        wait for Clk_period; 
        Features_din <= "0000000111001111";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000000100101010";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "1111110110011010";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000001011101010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000100100100011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000101001010101";
        wait for Clk_period; 
        Features_din <= "0000100010011110";
        wait for Clk_period; 
        Features_din <= "1111101100100111";
        wait for Clk_period; 
        Features_din <= "1111011110000110";
        wait for Clk_period; 
        Features_din <= "1111011010000000";
        wait for Clk_period; 
        Features_din <= "1111001101110101";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "1111011111010111";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000000110100000";
        wait for Clk_period; 
        Features_din <= "0000001011110011";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000010011000100";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000011011010";
        wait for Clk_period; 
        Features_din <= "1111110111100110";
        wait for Clk_period; 
        Features_din <= "0000000011011001";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001001111101";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000011010111";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001011100101000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "0000000111100100";
        wait for Clk_period; 
        Features_din <= "1111011100011111";
        wait for Clk_period; 
        Features_din <= "1111101000101100";
        wait for Clk_period; 
        Features_din <= "1111111000010111";
        wait for Clk_period; 
        Features_din <= "1111110010001100";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000100011011";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111100111101101";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "1111100101101111";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001111100101011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011110000001";
        wait for Clk_period; 
        Features_din <= "0000100011110001";
        wait for Clk_period; 
        Features_din <= "1111001000101010";
        wait for Clk_period; 
        Features_din <= "1111010011111101";
        wait for Clk_period; 
        Features_din <= "1111001010001000";
        wait for Clk_period; 
        Features_din <= "1111010001101101";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000110011101";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111101100100010";
        wait for Clk_period; 
        Features_din <= "1111100101101110";
        wait for Clk_period; 
        Features_din <= "0000001011101111";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001011101100";
        wait for Clk_period; 
        Features_din <= "0000001001000010";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000000011101011";
        wait for Clk_period; 
        Features_din <= "1111111100111000";
        wait for Clk_period; 
        Features_din <= "0000000101110100";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000000110000011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "0000000011011100";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000110001111010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000100000110111";
        wait for Clk_period; 
        Features_din <= "0000010100010101";
        wait for Clk_period; 
        Features_din <= "0000000110000010";
        wait for Clk_period; 
        Features_din <= "1111101101110010";
        wait for Clk_period; 
        Features_din <= "1111010010010010";
        wait for Clk_period; 
        Features_din <= "1111100111101000";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000001011110100";
        wait for Clk_period; 
        Features_din <= "1111011101000001";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "0000001000111011";
        wait for Clk_period; 
        Features_din <= "0000000111001011";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000000011110010";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "1111111000001100";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(3, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011100100111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111101110101100";
        wait for Clk_period; 
        Features_din <= "0000001011000111";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "0000011011100010";
        wait for Clk_period; 
        Features_din <= "1111111101111111";
        wait for Clk_period; 
        Features_din <= "1111011100110010";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111011110001010";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000000011110111";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000000101110111";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "1111110111010000";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000000111011100";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000011010110";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010110001110011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000100110000100";
        wait for Clk_period; 
        Features_din <= "1111111001010011";
        wait for Clk_period; 
        Features_din <= "1111010001000000";
        wait for Clk_period; 
        Features_din <= "1110110010101111";
        wait for Clk_period; 
        Features_din <= "1111110100100100";
        wait for Clk_period; 
        Features_din <= "1111101110011000";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111110011000111";
        wait for Clk_period; 
        Features_din <= "1111101011111111";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000000111011010";
        wait for Clk_period; 
        Features_din <= "1111101011100001";
        wait for Clk_period; 
        Features_din <= "0000010010010101";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000000101011001";
        wait for Clk_period; 
        Features_din <= "0000000011100100";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001100100100001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011000000100";
        wait for Clk_period; 
        Features_din <= "0000001000100010";
        wait for Clk_period; 
        Features_din <= "1111001100001110";
        wait for Clk_period; 
        Features_din <= "1111101110011111";
        wait for Clk_period; 
        Features_din <= "1111100001100010";
        wait for Clk_period; 
        Features_din <= "1111101011000100";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000001000101011";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111110000101101";
        wait for Clk_period; 
        Features_din <= "1111101010001111";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001100010001";
        wait for Clk_period; 
        Features_din <= "0000010101011111";
        wait for Clk_period; 
        Features_din <= "0000000101000000";
        wait for Clk_period; 
        Features_din <= "1111110100001001";
        wait for Clk_period; 
        Features_din <= "0000010100111111";
        wait for Clk_period; 
        Features_din <= "0000000110011110";
        wait for Clk_period; 
        Features_din <= "1111111111111111";
        wait for Clk_period; 
        Features_din <= "0000000101100000";
        wait for Clk_period; 
        Features_din <= "0000000010101101";
        wait for Clk_period; 
        Features_din <= "0000000111010111";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "0000000011111101";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001010101010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010001110100";
        wait for Clk_period; 
        Features_din <= "0000011010010011";
        wait for Clk_period; 
        Features_din <= "0000010010001001";
        wait for Clk_period; 
        Features_din <= "1111101011000110";
        wait for Clk_period; 
        Features_din <= "1111000111001011";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000001010100011";
        wait for Clk_period; 
        Features_din <= "1111011100011010";
        wait for Clk_period; 
        Features_din <= "0000001000111100";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000000101011100";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001000110101";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "1111111001000000";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000000011110011";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000011000101";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001110000000110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0001000010111001";
        wait for Clk_period; 
        Features_din <= "1111000111100011";
        wait for Clk_period; 
        Features_din <= "1111000101011001";
        wait for Clk_period; 
        Features_din <= "1111101110101101";
        wait for Clk_period; 
        Features_din <= "1110110011011101";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "1111111000110011";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111011111001101";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001001101101010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000101000011111";
        wait for Clk_period; 
        Features_din <= "0000111001000101";
        wait for Clk_period; 
        Features_din <= "1111011111101010";
        wait for Clk_period; 
        Features_din <= "1111100111111111";
        wait for Clk_period; 
        Features_din <= "1111101111000101";
        wait for Clk_period; 
        Features_din <= "1110111111101101";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000101010111";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000001000011011";
        wait for Clk_period; 
        Features_din <= "0000010100010001";
        wait for Clk_period; 
        Features_din <= "0000001010001101";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "1111110100011001";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000010100010111";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111100101100100";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "0000001100010010";
        wait for Clk_period; 
        Features_din <= "0000000101011001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "0000000011011110";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001010110001011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000100110010010";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "1111001111101000";
        wait for Clk_period; 
        Features_din <= "1110111101011101";
        wait for Clk_period; 
        Features_din <= "1111110000010101";
        wait for Clk_period; 
        Features_din <= "1111101101110101";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000111100110";
        wait for Clk_period; 
        Features_din <= "0000010011011111";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "1111111010101001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010100011111";
        wait for Clk_period; 
        Features_din <= "1111111000001110";
        wait for Clk_period; 
        Features_din <= "1111111010000011";
        wait for Clk_period; 
        Features_din <= "1111100011100010";
        wait for Clk_period; 
        Features_din <= "0000000100100010";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000001001000101";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001001111100111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001000100111100";
        wait for Clk_period; 
        Features_din <= "0000000011111111";
        wait for Clk_period; 
        Features_din <= "1111011001101111";
        wait for Clk_period; 
        Features_din <= "1111010101100000";
        wait for Clk_period; 
        Features_din <= "1111010010110101";
        wait for Clk_period; 
        Features_din <= "1111010000000001";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001011110010";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111101111111100";
        wait for Clk_period; 
        Features_din <= "0000000011010000";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "1111011111011100";
        wait for Clk_period; 
        Features_din <= "0000000011111101";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000001010010101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000011100011";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001100000110000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000000111000010";
        wait for Clk_period; 
        Features_din <= "0000001001111100";
        wait for Clk_period; 
        Features_din <= "1111101001111110";
        wait for Clk_period; 
        Features_din <= "1111011010110001";
        wait for Clk_period; 
        Features_din <= "1111110101111111";
        wait for Clk_period; 
        Features_din <= "1111001010010111";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000001011011000";
        wait for Clk_period; 
        Features_din <= "0000010001110100";
        wait for Clk_period; 
        Features_din <= "0000000100110110";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "1111110101110101";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "0000010001110100";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111111010010000";
        wait for Clk_period; 
        Features_din <= "1111100010001011";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001101000001011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001001110100000";
        wait for Clk_period; 
        Features_din <= "0000011001101010";
        wait for Clk_period; 
        Features_din <= "1111000111100110";
        wait for Clk_period; 
        Features_din <= "1111011100111011";
        wait for Clk_period; 
        Features_din <= "1111001011101011";
        wait for Clk_period; 
        Features_din <= "1111100010110010";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111011110101111";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000100000010";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000000100001110";
        wait for Clk_period; 
        Features_din <= "0000000011101110";
        wait for Clk_period; 
        Features_din <= "1111110110110100";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001100111110110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010010110011";
        wait for Clk_period; 
        Features_din <= "1111101101111011";
        wait for Clk_period; 
        Features_din <= "1111100111000000";
        wait for Clk_period; 
        Features_din <= "1111010111010101";
        wait for Clk_period; 
        Features_din <= "1111110000101001";
        wait for Clk_period; 
        Features_din <= "1111001101100011";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "1111101100100011";
        wait for Clk_period; 
        Features_din <= "0000010101001100";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000111000010";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "1111100101000000";
        wait for Clk_period; 
        Features_din <= "0000001010110000";
        wait for Clk_period; 
        Features_din <= "0000001000010111";
        wait for Clk_period; 
        Features_din <= "1111111111000111";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001001101000000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011100100110";
        wait for Clk_period; 
        Features_din <= "0000011000100100";
        wait for Clk_period; 
        Features_din <= "1111010011011110";
        wait for Clk_period; 
        Features_din <= "1111100011011001";
        wait for Clk_period; 
        Features_din <= "1111110001000010";
        wait for Clk_period; 
        Features_din <= "1111010001111011";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000100100111";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111101011101010";
        wait for Clk_period; 
        Features_din <= "0000010111010111";
        wait for Clk_period; 
        Features_din <= "0000001011110011";
        wait for Clk_period; 
        Features_din <= "0000000101111001";
        wait for Clk_period; 
        Features_din <= "0000000110101010";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111100110101000";
        wait for Clk_period; 
        Features_din <= "0000000111100011";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "1111111110111000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "0000001010110100";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001111001010000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000110010100101";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "1111011010001000";
        wait for Clk_period; 
        Features_din <= "1111001001011001";
        wait for Clk_period; 
        Features_din <= "1111101001010011";
        wait for Clk_period; 
        Features_din <= "1111011100010010";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000001001101000";
        wait for Clk_period; 
        Features_din <= "0000001001101000";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111110001001011";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000001001101000";
        wait for Clk_period; 
        Features_din <= "0000001001101000";
        wait for Clk_period; 
        Features_din <= "0000001001101000";
        wait for Clk_period; 
        Features_din <= "1111011110101101";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000011100010";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001000010000000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000110011101100";
        wait for Clk_period; 
        Features_din <= "0000010101001000";
        wait for Clk_period; 
        Features_din <= "1111100100000111";
        wait for Clk_period; 
        Features_din <= "1111101110111000";
        wait for Clk_period; 
        Features_din <= "1111100010110000";
        wait for Clk_period; 
        Features_din <= "1111100100011000";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "1111011111100010";
        wait for Clk_period; 
        Features_din <= "0000010001100100";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000001011111010";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000000101001001";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111110101110100";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001010011011";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000011000110";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010110010111101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000100110100101";
        wait for Clk_period; 
        Features_din <= "1110111110111100";
        wait for Clk_period; 
        Features_din <= "1111011011001010";
        wait for Clk_period; 
        Features_din <= "0000000111110110";
        wait for Clk_period; 
        Features_din <= "1111000111001111";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000011001001";
        wait for Clk_period; 
        Features_din <= "0000010110001101";
        wait for Clk_period; 
        Features_din <= "0000001010110001";
        wait for Clk_period; 
        Features_din <= "0000001001010111";
        wait for Clk_period; 
        Features_din <= "1111110111100110";
        wait for Clk_period; 
        Features_din <= "0000001011110110";
        wait for Clk_period; 
        Features_din <= "0000010010111000";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "1111111000001111";
        wait for Clk_period; 
        Features_din <= "1111100011101011";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "0000000011001100";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111011000011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010110110";
        wait for Clk_period; 
        Features_din <= "1111111000101011";
        wait for Clk_period; 
        Features_din <= "0000010101111100";
        wait for Clk_period; 
        Features_din <= "0000011000110001";
        wait for Clk_period; 
        Features_din <= "1111100111101011";
        wait for Clk_period; 
        Features_din <= "1111010100101101";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "0000001001010110";
        wait for Clk_period; 
        Features_din <= "1111111011101111";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "1111110111100000";
        wait for Clk_period; 
        Features_din <= "1111111100000000";
        wait for Clk_period; 
        Features_din <= "1111100001011110";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000011010000";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010011000110110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000000100001001";
        wait for Clk_period; 
        Features_din <= "0000000111110111";
        wait for Clk_period; 
        Features_din <= "1110111000010001";
        wait for Clk_period; 
        Features_din <= "1111011000111101";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "1111010101101110";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111110001101101";
        wait for Clk_period; 
        Features_din <= "1111101111001010";
        wait for Clk_period; 
        Features_din <= "0000001001100011";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000010001111100";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "1111101001111111";
        wait for Clk_period; 
        Features_din <= "0000001000110100";
        wait for Clk_period; 
        Features_din <= "0000010011001010";
        wait for Clk_period; 
        Features_din <= "0000000111010010";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001010110001111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011001100011";
        wait for Clk_period; 
        Features_din <= "0000011001000011";
        wait for Clk_period; 
        Features_din <= "1111011101111000";
        wait for Clk_period; 
        Features_din <= "1111011010111010";
        wait for Clk_period; 
        Features_din <= "1111110010001101";
        wait for Clk_period; 
        Features_din <= "1111011110010011";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000001010110000";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111110000111010";
        wait for Clk_period; 
        Features_din <= "1111101001001001";
        wait for Clk_period; 
        Features_din <= "0000000110111010";
        wait for Clk_period; 
        Features_din <= "0000000011101111";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000000100101001";
        wait for Clk_period; 
        Features_din <= "1111110000001101";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000000110010111";
        wait for Clk_period; 
        Features_din <= "0000000101011100";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001001110110";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000011001001";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001111101001000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010101101110";
        wait for Clk_period; 
        Features_din <= "0000000110010100";
        wait for Clk_period; 
        Features_din <= "1111001110101101";
        wait for Clk_period; 
        Features_din <= "1111001101111011";
        wait for Clk_period; 
        Features_din <= "0000000011011000";
        wait for Clk_period; 
        Features_din <= "1111011000110011";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000110111100";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111101101001111";
        wait for Clk_period; 
        Features_din <= "0000010111100101";
        wait for Clk_period; 
        Features_din <= "0000000111101010";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000001001010000";
        wait for Clk_period; 
        Features_din <= "1111101000101110";
        wait for Clk_period; 
        Features_din <= "1111111010000010";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001000011101";
        wait for Clk_period; 
        Features_din <= "0000001001100000";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000001010100101";
        wait for Clk_period; 
        Features_din <= "0000000100010000";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010001111001101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010011110001";
        wait for Clk_period; 
        Features_din <= "1111101101011011";
        wait for Clk_period; 
        Features_din <= "1111001011011001";
        wait for Clk_period; 
        Features_din <= "1111011111110011";
        wait for Clk_period; 
        Features_din <= "1111110000110111";
        wait for Clk_period; 
        Features_din <= "1111001111010110";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000011100000";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "1111100100000010";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "1111101001100110";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000011100001";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001101110010101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111101110010001";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "1111001111111101";
        wait for Clk_period; 
        Features_din <= "1111011001001011";
        wait for Clk_period; 
        Features_din <= "1111111101011010";
        wait for Clk_period; 
        Features_din <= "1111110010110101";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000100110001";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111101101100010";
        wait for Clk_period; 
        Features_din <= "1111100100100111";
        wait for Clk_period; 
        Features_din <= "0000000101010110";
        wait for Clk_period; 
        Features_din <= "0000001000001010";
        wait for Clk_period; 
        Features_din <= "0000000101010110";
        wait for Clk_period; 
        Features_din <= "0000000111100100";
        wait for Clk_period; 
        Features_din <= "0000010101110100";
        wait for Clk_period; 
        Features_din <= "0000001010110100";
        wait for Clk_period; 
        Features_din <= "0000001000111001";
        wait for Clk_period; 
        Features_din <= "1111111111000000";
        wait for Clk_period; 
        Features_din <= "0000000110010000";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001011010011";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000011010111";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000010010010110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010110111100";
        wait for Clk_period; 
        Features_din <= "0000010011100101";
        wait for Clk_period; 
        Features_din <= "1111110011011100";
        wait for Clk_period; 
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "1111111010100100";
        wait for Clk_period; 
        Features_din <= "1111100010000011";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111101011101001";
        wait for Clk_period; 
        Features_din <= "1111100101011100";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000001100100010";
        wait for Clk_period; 
        Features_din <= "0000001000111101";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000010100101001";
        wait for Clk_period; 
        Features_din <= "0000001001011000";
        wait for Clk_period; 
        Features_din <= "0000001000110010";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "0000001001010101";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000000011011100";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011000111001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000111010011000";
        wait for Clk_period; 
        Features_din <= "0000100111100010";
        wait for Clk_period; 
        Features_din <= "1111110001011101";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "1111100000100100";
        wait for Clk_period; 
        Features_din <= "1111001000101010";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000111011110";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "1111110011001110";
        wait for Clk_period; 
        Features_din <= "1111101100110100";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001010111011";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "1111101010010111";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000000110000010";
        wait for Clk_period; 
        Features_din <= "0000001001000000";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000011010001";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001011001100000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011010101000";
        wait for Clk_period; 
        Features_din <= "0000011000110100";
        wait for Clk_period; 
        Features_din <= "1111001111111001";
        wait for Clk_period; 
        Features_din <= "1111001111011011";
        wait for Clk_period; 
        Features_din <= "1111111000111000";
        wait for Clk_period; 
        Features_din <= "1111010100011110";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111101101111011";
        wait for Clk_period; 
        Features_din <= "1111100100111101";
        wait for Clk_period; 
        Features_din <= "0000000110111100";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "0000001001110100";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000010100010001";
        wait for Clk_period; 
        Features_din <= "0000001100001000";
        wait for Clk_period; 
        Features_din <= "0000000111101000";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001000001001";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000011011001";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001110001011111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011010100000";
        wait for Clk_period; 
        Features_din <= "0000000101011010";
        wait for Clk_period; 
        Features_din <= "1111110010111011";
        wait for Clk_period; 
        Features_din <= "1111001100110100";
        wait for Clk_period; 
        Features_din <= "1111010001110000";
        wait for Clk_period; 
        Features_din <= "1111100010001000";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111101010110101";
        wait for Clk_period; 
        Features_din <= "0000010100011000";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000001010100011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111100110001100";
        wait for Clk_period; 
        Features_din <= "0000001001001101";
        wait for Clk_period; 
        Features_din <= "0000001000000001";
        wait for Clk_period; 
        Features_din <= "1111111110110101";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001111111101111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111110110000010";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "1111000010100101";
        wait for Clk_period; 
        Features_din <= "1111000110000001";
        wait for Clk_period; 
        Features_din <= "1111110111000101";
        wait for Clk_period; 
        Features_din <= "1111100001000000";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "1111110011100001";
        wait for Clk_period; 
        Features_din <= "1111101100110101";
        wait for Clk_period; 
        Features_din <= "0000000101000001";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "1111101001111001";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000000111010011";
        wait for Clk_period; 
        Features_din <= "0000000110011001";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001001010000000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011111111001";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "1111010110100010";
        wait for Clk_period; 
        Features_din <= "1111100100111101";
        wait for Clk_period; 
        Features_din <= "1111101101011111";
        wait for Clk_period; 
        Features_din <= "1111011011100000";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "1111101101100111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111000101111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000011011110010";
        wait for Clk_period; 
        Features_din <= "1111101111001111";
        wait for Clk_period; 
        Features_din <= "1111111001100111";
        wait for Clk_period; 
        Features_din <= "0000000011111101";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010000011000000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111110100000100";
        wait for Clk_period; 
        Features_din <= "0000000100010001";
        wait for Clk_period; 
        Features_din <= "1111010010111000";
        wait for Clk_period; 
        Features_din <= "1111100101000010";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "1111100011100111";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111011110110001";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000000010111101";
        wait for Clk_period; 
        Features_din <= "0000000011011011";
        wait for Clk_period; 
        Features_din <= "0000000011001010";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000000100011011";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "1111110110100100";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000011010110";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001010011100000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001001101100101";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "1111011001000101";
        wait for Clk_period; 
        Features_din <= "1111011110111000";
        wait for Clk_period; 
        Features_din <= "1111011011100001";
        wait for Clk_period; 
        Features_din <= "1111010001101111";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111111101001011";
        wait for Clk_period; 
        Features_din <= "1111101010011110";
        wait for Clk_period; 
        Features_din <= "0000001100000001";
        wait for Clk_period; 
        Features_din <= "0000000110010101";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000000101000100";
        wait for Clk_period; 
        Features_din <= "1111101000101110";
        wait for Clk_period; 
        Features_din <= "0000000110101001";
        wait for Clk_period; 
        Features_din <= "0000000011011101";
        wait for Clk_period; 
        Features_din <= "0000010101101101";
        wait for Clk_period; 
        Features_din <= "0000000101001100";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000011000110";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001100111110100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100101010";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "1111010111110101";
        wait for Clk_period; 
        Features_din <= "1111100110110000";
        wait for Clk_period; 
        Features_din <= "1111110001110110";
        wait for Clk_period; 
        Features_din <= "1111011011010001";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000111111001";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111101100000011";
        wait for Clk_period; 
        Features_din <= "1111100110001011";
        wait for Clk_period; 
        Features_din <= "0000000100100010";
        wait for Clk_period; 
        Features_din <= "0000001011101100";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000010101010010";
        wait for Clk_period; 
        Features_din <= "0000001011111001";
        wait for Clk_period; 
        Features_din <= "0000000101111011";
        wait for Clk_period; 
        Features_din <= "1111111101001110";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000000111010011";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000011011101";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001100111000101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011000100101";
        wait for Clk_period; 
        Features_din <= "0000000101010111";
        wait for Clk_period; 
        Features_din <= "1111001100100111";
        wait for Clk_period; 
        Features_din <= "1111011111011010";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "1111011011010001";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000001001000000";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111101100100111";
        wait for Clk_period; 
        Features_din <= "1111100101110010";
        wait for Clk_period; 
        Features_din <= "0000000111001010";
        wait for Clk_period; 
        Features_din <= "0000000011001010";
        wait for Clk_period; 
        Features_din <= "0000000110001100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010111011001";
        wait for Clk_period; 
        Features_din <= "0000000111111111";
        wait for Clk_period; 
        Features_din <= "0000001000110110";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001100100110";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000011011100";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(2, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111001011101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010110010";
        wait for Clk_period; 
        Features_din <= "0000000100000101";
        wait for Clk_period; 
        Features_din <= "0000100110001011";
        wait for Clk_period; 
        Features_din <= "0000000111100010";
        wait for Clk_period; 
        Features_din <= "1111110010010101";
        wait for Clk_period; 
        Features_din <= "1111101111111010";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000100101010";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111110100001101";
        wait for Clk_period; 
        Features_din <= "1111101100001010";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001100011100";
        wait for Clk_period; 
        Features_din <= "0000000110011100";
        wait for Clk_period; 
        Features_din <= "1111101010010011";
        wait for Clk_period; 
        Features_din <= "0000010001100011";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000000110100011";
        wait for Clk_period; 
        Features_din <= "0000001011100000";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000010101101";
        wait for Clk_period; 
        Features_din <= "0000000100000111";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(3, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000010010101010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000000100000000";
        wait for Clk_period; 
        Features_din <= "0000110001001000";
        wait for Clk_period; 
        Features_din <= "1111101111110100";
        wait for Clk_period; 
        Features_din <= "0000011000101110";
        wait for Clk_period; 
        Features_din <= "1111100101110001";
        wait for Clk_period; 
        Features_din <= "1111000110111111";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000110110010";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "1111101001001101";
        wait for Clk_period; 
        Features_din <= "1111101000000011";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001100000011";
        wait for Clk_period; 
        Features_din <= "0000001000100101";
        wait for Clk_period; 
        Features_din <= "0000000011010000";
        wait for Clk_period; 
        Features_din <= "0000010101011110";
        wait for Clk_period; 
        Features_din <= "0000001001111001";
        wait for Clk_period; 
        Features_din <= "0000001000000100";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "0000001000000100";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "0000000011110111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "0000000100011001";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010110010111001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000100100110111";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "1111100000111010";
        wait for Clk_period; 
        Features_din <= "1111011101100100";
        wait for Clk_period; 
        Features_din <= "1111101101111110";
        wait for Clk_period; 
        Features_din <= "1111010010110001";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "1111100111011011";
        wait for Clk_period; 
        Features_din <= "0000000101000110";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "1111101000101000";
        wait for Clk_period; 
        Features_din <= "0000001001110011";
        wait for Clk_period; 
        Features_din <= "0000001000001001";
        wait for Clk_period; 
        Features_din <= "1111111111001100";
        wait for Clk_period; 
        Features_din <= "0000000101101100";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000110101001111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011111010001";
        wait for Clk_period; 
        Features_din <= "0000010001011010";
        wait for Clk_period; 
        Features_din <= "1111100100001111";
        wait for Clk_period; 
        Features_din <= "1111001010010010";
        wait for Clk_period; 
        Features_din <= "1111110010100000";
        wait for Clk_period; 
        Features_din <= "1111011110011111";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "1111110101101110";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1111100001010001";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000000110111011";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001010001100101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111101101111011";
        wait for Clk_period; 
        Features_din <= "0000000101101011";
        wait for Clk_period; 
        Features_din <= "1111011111011110";
        wait for Clk_period; 
        Features_din <= "1111011100111011";
        wait for Clk_period; 
        Features_din <= "0000010100110001";
        wait for Clk_period; 
        Features_din <= "1111101101010000";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111110001100100";
        wait for Clk_period; 
        Features_din <= "1111101011100000";
        wait for Clk_period; 
        Features_din <= "0000000011101110";
        wait for Clk_period; 
        Features_din <= "0000000011111011";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000000100011110";
        wait for Clk_period; 
        Features_din <= "1111101101000011";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000000101111110";
        wait for Clk_period; 
        Features_din <= "0000001001111011";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001011111011";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(3, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111110111011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "1111110101111001";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000100010011010";
        wait for Clk_period; 
        Features_din <= "1111101100110000";
        wait for Clk_period; 
        Features_din <= "1111001100100000";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000101010100";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000000111010000";
        wait for Clk_period; 
        Features_din <= "0000000111111100";
        wait for Clk_period; 
        Features_din <= "1111110010000110";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000010100101101";
        wait for Clk_period; 
        Features_din <= "1111110101101100";
        wait for Clk_period; 
        Features_din <= "1111111011110001";
        wait for Clk_period; 
        Features_din <= "1111101000100100";
        wait for Clk_period; 
        Features_din <= "0000001010101010";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000001010100101";
        wait for Clk_period; 
        Features_din <= "0000000111001010";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001010110100000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001000001000000";
        wait for Clk_period; 
        Features_din <= "1111110110100110";
        wait for Clk_period; 
        Features_din <= "1111011110001101";
        wait for Clk_period; 
        Features_din <= "1111011110100001";
        wait for Clk_period; 
        Features_din <= "1111011111011101";
        wait for Clk_period; 
        Features_din <= "1110110111011101";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000110011110";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "1111101100011011";
        wait for Clk_period; 
        Features_din <= "1111100100101100";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "0000000011111111";
        wait for Clk_period; 
        Features_din <= "0000000111101011";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000010100111011";
        wait for Clk_period; 
        Features_din <= "0000001000011010";
        wait for Clk_period; 
        Features_din <= "0000001001110000";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000011011111";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000111111011001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010111101011";
        wait for Clk_period; 
        Features_din <= "0000000110110011";
        wait for Clk_period; 
        Features_din <= "1111101100111100";
        wait for Clk_period; 
        Features_din <= "1111111010010101";
        wait for Clk_period; 
        Features_din <= "1111110111111111";
        wait for Clk_period; 
        Features_din <= "1111100010100010";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000110000000";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111101100100000";
        wait for Clk_period; 
        Features_din <= "1111100100111001";
        wait for Clk_period; 
        Features_din <= "0000001100001110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001000000001";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000010100110000";
        wait for Clk_period; 
        Features_din <= "0000001010100111";
        wait for Clk_period; 
        Features_din <= "0000001000010000";
        wait for Clk_period; 
        Features_din <= "1111111110111111";
        wait for Clk_period; 
        Features_din <= "0000000011110111";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "0000001010001111";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "0000000011101001";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000101010000001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011100111001";
        wait for Clk_period; 
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "1111110001110001";
        wait for Clk_period; 
        Features_din <= "1110110001101101";
        wait for Clk_period; 
        Features_din <= "1111011011000110";
        wait for Clk_period; 
        Features_din <= "0001000000010100";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000010111111";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111011110111110";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000000100010000";
        wait for Clk_period; 
        Features_din <= "0000001011000110";
        wait for Clk_period; 
        Features_din <= "0000000011101100";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000000101110011";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "1111110101111111";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001011000110";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001110101001010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001000000001000";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "1110111110000000";
        wait for Clk_period; 
        Features_din <= "1111100010010001";
        wait for Clk_period; 
        Features_din <= "1111100110011001";
        wait for Clk_period; 
        Features_din <= "1110111101111101";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000001011011000";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "1111101011101001";
        wait for Clk_period; 
        Features_din <= "1111100110111001";
        wait for Clk_period; 
        Features_din <= "0000000110111111";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000010011000000";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000000100100010";
        wait for Clk_period; 
        Features_din <= "1111111011101001";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000000100010001";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000011010011";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011001110110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011010010101";
        wait for Clk_period; 
        Features_din <= "0000000100011100";
        wait for Clk_period; 
        Features_din <= "1111110010010010";
        wait for Clk_period; 
        Features_din <= "0000011101011000";
        wait for Clk_period; 
        Features_din <= "1111100100000010";
        wait for Clk_period; 
        Features_din <= "1111001101101111";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000001011000100";
        wait for Clk_period; 
        Features_din <= "0000010011001011";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "0000000101000101";
        wait for Clk_period; 
        Features_din <= "1111110010010111";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000010011001011";
        wait for Clk_period; 
        Features_din <= "1111110100110010";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111100111000011";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000011010110";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001010011101111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000111001100011";
        wait for Clk_period; 
        Features_din <= "0000000100001101";
        wait for Clk_period; 
        Features_din <= "1111011010101100";
        wait for Clk_period; 
        Features_din <= "1111100100000110";
        wait for Clk_period; 
        Features_din <= "1111101001110101";
        wait for Clk_period; 
        Features_din <= "1110111111100101";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000011100010";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000001011001001";
        wait for Clk_period; 
        Features_din <= "0000010001001101";
        wait for Clk_period; 
        Features_din <= "0000001010001011";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000000100101111";
        wait for Clk_period; 
        Features_din <= "0000000101000011";
        wait for Clk_period; 
        Features_din <= "1111011100101100";
        wait for Clk_period; 
        Features_din <= "0000000110011000";
        wait for Clk_period; 
        Features_din <= "0000000011000101";
        wait for Clk_period; 
        Features_din <= "1111111000110001";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000001011010010";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000011010010";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000100001010010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001000011101000";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "1111110110101100";
        wait for Clk_period; 
        Features_din <= "1111100011011110";
        wait for Clk_period; 
        Features_din <= "1111101001110111";
        wait for Clk_period; 
        Features_din <= "1111001101010000";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111011110010101";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000000100110001";
        wait for Clk_period; 
        Features_din <= "0000000011101011";
        wait for Clk_period; 
        Features_din <= "1111110110100010";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000001001001000";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001010110101000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001000000100111";
        wait for Clk_period; 
        Features_din <= "1111110010011101";
        wait for Clk_period; 
        Features_din <= "1111001001100100";
        wait for Clk_period; 
        Features_din <= "0000000100101000";
        wait for Clk_period; 
        Features_din <= "1111011000100001";
        wait for Clk_period; 
        Features_din <= "1111001010011010";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000001010111001";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "0000000010111101";
        wait for Clk_period; 
        Features_din <= "0000001010110110";
        wait for Clk_period; 
        Features_din <= "0000001010101101";
        wait for Clk_period; 
        Features_din <= "1111011100000100";
        wait for Clk_period; 
        Features_din <= "0000000110011110";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "1111111001010101";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000001011011011";
        wait for Clk_period; 
        Features_din <= "0000001000001110";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "0000000011001000";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001100010110000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "1111100110111111";
        wait for Clk_period; 
        Features_din <= "1111100110101101";
        wait for Clk_period; 
        Features_din <= "1111101100000100";
        wait for Clk_period; 
        Features_din <= "1111110010101011";
        wait for Clk_period; 
        Features_din <= "1111100110100011";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000101101110";
        wait for Clk_period; 
        Features_din <= "0000010100000000";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "1111111001011000";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "0000010100111001";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "1111111000100001";
        wait for Clk_period; 
        Features_din <= "1111100011100111";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000000011100101";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001111011000010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000111111001011";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "1111001110110000";
        wait for Clk_period; 
        Features_din <= "1111010110111000";
        wait for Clk_period; 
        Features_din <= "1111100001100100";
        wait for Clk_period; 
        Features_din <= "1111000100111101";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000001000110111";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111110011000100";
        wait for Clk_period; 
        Features_din <= "1111101011010011";
        wait for Clk_period; 
        Features_din <= "0000000011101110";
        wait for Clk_period; 
        Features_din <= "0000000111001011";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "1111101100010101";
        wait for Clk_period; 
        Features_din <= "0000010010111011";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000000101010101";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001011001010";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000011101110";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000110010010001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000101100011000";
        wait for Clk_period; 
        Features_din <= "0001001010001110";
        wait for Clk_period; 
        Features_din <= "1111000110111011";
        wait for Clk_period; 
        Features_din <= "1111100011101001";
        wait for Clk_period; 
        Features_din <= "1111011100110100";
        wait for Clk_period; 
        Features_din <= "1111000110111101";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000001011011001";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111110100010011";
        wait for Clk_period; 
        Features_din <= "1111101100011011";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000000011001100";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101010000011";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010010100001";
        wait for Clk_period; 
        Features_din <= "0000000110010001";
        wait for Clk_period; 
        Features_din <= "0000001010110001";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "0000000011011110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010000000011100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000110100000000";
        wait for Clk_period; 
        Features_din <= "1111010110101100";
        wait for Clk_period; 
        Features_din <= "1111100000111001";
        wait for Clk_period; 
        Features_din <= "1111110011000001";
        wait for Clk_period; 
        Features_din <= "1111000011000110";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000111100101";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111110011001110";
        wait for Clk_period; 
        Features_din <= "1111101101000001";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101010011011";
        wait for Clk_period; 
        Features_din <= "0000010010000100";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000000101011101";
        wait for Clk_period; 
        Features_din <= "0000000101001010";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "0000000111111010";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000101000010011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000100001110000";
        wait for Clk_period; 
        Features_din <= "0000110100111111";
        wait for Clk_period; 
        Features_din <= "1111110111001100";
        wait for Clk_period; 
        Features_din <= "1111110001001101";
        wait for Clk_period; 
        Features_din <= "1111110111000100";
        wait for Clk_period; 
        Features_din <= "1110111111100110";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000100101000";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "1111110011001011";
        wait for Clk_period; 
        Features_din <= "1111101100001011";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001011100101";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000000111101001";
        wait for Clk_period; 
        Features_din <= "1111101010111011";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000000110100111";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010001010010000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111110111110101";
        wait for Clk_period; 
        Features_din <= "1111110100010000";
        wait for Clk_period; 
        Features_din <= "1110111010111110";
        wait for Clk_period; 
        Features_din <= "1111010100000100";
        wait for Clk_period; 
        Features_din <= "1111101110110101";
        wait for Clk_period; 
        Features_din <= "1111001101100011";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000101110011";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111100101011011";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "1111101000000010";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000011001101";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000110110111011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011101011111";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "1111100000010011";
        wait for Clk_period; 
        Features_din <= "1111101101101110";
        wait for Clk_period; 
        Features_din <= "1111101010011010";
        wait for Clk_period; 
        Features_din <= "1111100111111111";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000111111111";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000001010011110";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000000111111110";
        wait for Clk_period; 
        Features_din <= "0000000011000010";
        wait for Clk_period; 
        Features_din <= "0000000111100111";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "1111011011001110";
        wait for Clk_period; 
        Features_din <= "0000001000000010";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "1111111011000001";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000011010111";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001110101100111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010100000111";
        wait for Clk_period; 
        Features_din <= "0000000011000111";
        wait for Clk_period; 
        Features_din <= "1111011001000010";
        wait for Clk_period; 
        Features_din <= "1111101011011000";
        wait for Clk_period; 
        Features_din <= "1111101100100101";
        wait for Clk_period; 
        Features_din <= "1111001100000011";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000011101111";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111011110001111";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000000100101111";
        wait for Clk_period; 
        Features_din <= "0000001011110010";
        wait for Clk_period; 
        Features_din <= "0000000110011000";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000000100011100";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111110110011100";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010100000110011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001011100011";
        wait for Clk_period; 
        Features_din <= "0000101000000000";
        wait for Clk_period; 
        Features_din <= "1111000111000011";
        wait for Clk_period; 
        Features_din <= "1110101110111010";
        wait for Clk_period; 
        Features_din <= "1111100110101001";
        wait for Clk_period; 
        Features_din <= "1111010000011010";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000111110001";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000010001110001";
        wait for Clk_period; 
        Features_din <= "0000011100011100";
        wait for Clk_period; 
        Features_din <= "0000001011101011";
        wait for Clk_period; 
        Features_din <= "0000001001110011";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "1111101100101000";
        wait for Clk_period; 
        Features_din <= "1111110010101110";
        wait for Clk_period; 
        Features_din <= "1111110110000001";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000001001111111";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000101000010";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000011011011";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001011111111110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000100110101001";
        wait for Clk_period; 
        Features_din <= "0000101000101111";
        wait for Clk_period; 
        Features_din <= "1111011000010111";
        wait for Clk_period; 
        Features_din <= "1111010001100001";
        wait for Clk_period; 
        Features_din <= "1111100011001100";
        wait for Clk_period; 
        Features_din <= "1111011011111001";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000110110110";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111110011100001";
        wait for Clk_period; 
        Features_din <= "1111101011111111";
        wait for Clk_period; 
        Features_din <= "0000000011000010";
        wait for Clk_period; 
        Features_din <= "0000001010101110";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101011000100";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000000101110101";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "0000000011110111";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001010001001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000110101010000";
        wait for Clk_period; 
        Features_din <= "1111111101010001";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "1111111101011000";
        wait for Clk_period; 
        Features_din <= "1111110100101110";
        wait for Clk_period; 
        Features_din <= "1111010000111011";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000011110000001";
        wait for Clk_period; 
        Features_din <= "1111101100100010";
        wait for Clk_period; 
        Features_din <= "0000001000111111";
        wait for Clk_period; 
        Features_din <= "0000000011011110";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000001100100011";
        wait for Clk_period; 
        Features_din <= "1111101111111000";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001000101011";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "0000000100010000";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000011100010";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001001111010011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000110011110100";
        wait for Clk_period; 
        Features_din <= "0000000011110110";
        wait for Clk_period; 
        Features_din <= "1111011001010011";
        wait for Clk_period; 
        Features_din <= "1111101111010110";
        wait for Clk_period; 
        Features_din <= "1111110011101100";
        wait for Clk_period; 
        Features_din <= "1111100100000010";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000001001000100";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000001000000111";
        wait for Clk_period; 
        Features_din <= "0000010010110110";
        wait for Clk_period; 
        Features_din <= "0000000110100100";
        wait for Clk_period; 
        Features_din <= "0000000010111111";
        wait for Clk_period; 
        Features_din <= "0000000110101001";
        wait for Clk_period; 
        Features_din <= "0000000101000010";
        wait for Clk_period; 
        Features_din <= "1111011110010100";
        wait for Clk_period; 
        Features_din <= "0000001010010011";
        wait for Clk_period; 
        Features_din <= "1111111111000001";
        wait for Clk_period; 
        Features_din <= "1111110110110010";
        wait for Clk_period; 
        Features_din <= "0000000101011001";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001011101010";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "0000000010111110";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001111010101110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001000110111";
        wait for Clk_period; 
        Features_din <= "0000000100111100";
        wait for Clk_period; 
        Features_din <= "1110111100011100";
        wait for Clk_period; 
        Features_din <= "1111100100011100";
        wait for Clk_period; 
        Features_din <= "1111110001010110";
        wait for Clk_period; 
        Features_din <= "1111001000000110";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000010101100";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "1111101001001011";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "1111100100011001";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001110000010101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010011110011";
        wait for Clk_period; 
        Features_din <= "1111111100100011";
        wait for Clk_period; 
        Features_din <= "1111011010010010";
        wait for Clk_period; 
        Features_din <= "1111101001011111";
        wait for Clk_period; 
        Features_din <= "1111100010001010";
        wait for Clk_period; 
        Features_din <= "1111100110010101";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000011101101";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000010101101010";
        wait for Clk_period; 
        Features_din <= "1111111101100001";
        wait for Clk_period; 
        Features_din <= "0000000110110000";
        wait for Clk_period; 
        Features_din <= "0000000110000011";
        wait for Clk_period; 
        Features_din <= "0000001000111100";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "1111100010010100";
        wait for Clk_period; 
        Features_din <= "1111111011110100";
        wait for Clk_period; 
        Features_din <= "1111110110001110";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000011000010";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001111011000111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "1111000101011110";
        wait for Clk_period; 
        Features_din <= "1111100010100000";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "1111110000010111";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000101000110";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111110010110100";
        wait for Clk_period; 
        Features_din <= "1111101010011100";
        wait for Clk_period; 
        Features_din <= "0000000110110000";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000000110100111";
        wait for Clk_period; 
        Features_din <= "1111101100101111";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000000111010000";
        wait for Clk_period; 
        Features_din <= "0000000110000001";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001110100110010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001000010110011";
        wait for Clk_period; 
        Features_din <= "1111111100110011";
        wait for Clk_period; 
        Features_din <= "1110111101011000";
        wait for Clk_period; 
        Features_din <= "1111000011001100";
        wait for Clk_period; 
        Features_din <= "1111010100011100";
        wait for Clk_period; 
        Features_din <= "1111101001101110";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "1111100110100001";
        wait for Clk_period; 
        Features_din <= "0000000011010000";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001010011011";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "1111101000110001";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000001001010010";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000011101111";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000000100100011";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010000011001111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000101010110100";
        wait for Clk_period; 
        Features_din <= "0000010011111010";
        wait for Clk_period; 
        Features_din <= "1110111111000101";
        wait for Clk_period; 
        Features_din <= "1111001011100000";
        wait for Clk_period; 
        Features_din <= "1111101010010001";
        wait for Clk_period; 
        Features_din <= "1111011011111111";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000011111100";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "1111101100100110";
        wait for Clk_period; 
        Features_din <= "1111100110000111";
        wait for Clk_period; 
        Features_din <= "0000000011111011";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000000110111100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010111011100";
        wait for Clk_period; 
        Features_din <= "0000001001001101";
        wait for Clk_period; 
        Features_din <= "0000000111101011";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000011011110";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000100000100000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011000011010";
        wait for Clk_period; 
        Features_din <= "0001000100111011";
        wait for Clk_period; 
        Features_din <= "1111101100101101";
        wait for Clk_period; 
        Features_din <= "1111111110000111";
        wait for Clk_period; 
        Features_din <= "1111110100110010";
        wait for Clk_period; 
        Features_din <= "1111001110110011";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000100001010";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000001010111010";
        wait for Clk_period; 
        Features_din <= "1111011101101111";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000010100010101";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000000110010100";
        wait for Clk_period; 
        Features_din <= "1111111001101000";
        wait for Clk_period; 
        Features_din <= "0000001001000100";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000101011001";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111100001111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000101100101101";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "1111101100100101";
        wait for Clk_period; 
        Features_din <= "0000011101100000";
        wait for Clk_period; 
        Features_din <= "1111101010111010";
        wait for Clk_period; 
        Features_din <= "1111001110101111";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000010101001010";
        wait for Clk_period; 
        Features_din <= "1111110001010010";
        wait for Clk_period; 
        Features_din <= "0000001100111000";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "1111111010101010";
        wait for Clk_period; 
        Features_din <= "0000001000100011";
        wait for Clk_period; 
        Features_din <= "0000001100111000";
        wait for Clk_period; 
        Features_din <= "1111100100001010";
        wait for Clk_period; 
        Features_din <= "0000001100100000";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000001001011101";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "0000000100001000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "0000000100010000";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001100111001100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000100100011101";
        wait for Clk_period; 
        Features_din <= "0000011001110100";
        wait for Clk_period; 
        Features_din <= "1111101110010011";
        wait for Clk_period; 
        Features_din <= "1111010001001000";
        wait for Clk_period; 
        Features_din <= "1111011110100001";
        wait for Clk_period; 
        Features_din <= "1111001010010000";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000001000100010";
        wait for Clk_period; 
        Features_din <= "0000010011001011";
        wait for Clk_period; 
        Features_din <= "0000000100001111";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "1111111000111100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010011001011";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "1111111010000100";
        wait for Clk_period; 
        Features_din <= "1111100010010100";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010001010100000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "1111101100010011";
        wait for Clk_period; 
        Features_din <= "1110111011000001";
        wait for Clk_period; 
        Features_din <= "1111100101011011";
        wait for Clk_period; 
        Features_din <= "1111110111000110";
        wait for Clk_period; 
        Features_din <= "1111010100101001";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111101101101110";
        wait for Clk_period; 
        Features_din <= "1111100011001010";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "0000001011001010";
        wait for Clk_period; 
        Features_din <= "0000000101001100";
        wait for Clk_period; 
        Features_din <= "0000010001110010";
        wait for Clk_period; 
        Features_din <= "0000001011101100";
        wait for Clk_period; 
        Features_din <= "0000000110111101";
        wait for Clk_period; 
        Features_din <= "1111111111100011";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010001010000100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111101000101011";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "1111010010000101";
        wait for Clk_period; 
        Features_din <= "1110111100111011";
        wait for Clk_period; 
        Features_din <= "1111110100001011";
        wait for Clk_period; 
        Features_din <= "1111011011101000";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111101011101111";
        wait for Clk_period; 
        Features_din <= "1111100101100111";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "0000000111010100";
        wait for Clk_period; 
        Features_din <= "0000001000111101";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000010100111001";
        wait for Clk_period; 
        Features_din <= "0000001010011001";
        wait for Clk_period; 
        Features_din <= "0000000111101101";
        wait for Clk_period; 
        Features_din <= "1111111110101110";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001110010010011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111001011000";
        wait for Clk_period; 
        Features_din <= "1111011010011110";
        wait for Clk_period; 
        Features_din <= "1111001000110001";
        wait for Clk_period; 
        Features_din <= "1111011111110010";
        wait for Clk_period; 
        Features_din <= "1111111111011010";
        wait for Clk_period; 
        Features_din <= "1111101011100001";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000011101101110";
        wait for Clk_period; 
        Features_din <= "1111101100011110";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "1111101111101010";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "1111111011100100";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "0000000011001101";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001111101111111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000000101000101";
        wait for Clk_period; 
        Features_din <= "1111000001010011";
        wait for Clk_period; 
        Features_din <= "1111001110001000";
        wait for Clk_period; 
        Features_din <= "1111110101110001";
        wait for Clk_period; 
        Features_din <= "1111001011111101";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111011111110111";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001010101010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "0000000100101101";
        wait for Clk_period; 
        Features_din <= "0000010001111100";
        wait for Clk_period; 
        Features_din <= "0000001000101111";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111110100111010";
        wait for Clk_period; 
        Features_din <= "0000000100011001";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000001010111110";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000011010000";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010010010111010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011001110010";
        wait for Clk_period; 
        Features_din <= "1111110011011111";
        wait for Clk_period; 
        Features_din <= "1111010100110100";
        wait for Clk_period; 
        Features_din <= "1111010100010011";
        wait for Clk_period; 
        Features_din <= "1111100111101000";
        wait for Clk_period; 
        Features_din <= "1111101010110010";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000100001000";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "1111101010111110";
        wait for Clk_period; 
        Features_din <= "1111100111100011";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000000110100011";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000000101110000";
        wait for Clk_period; 
        Features_din <= "0000010010101000";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "1111111100010101";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010010001010110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000000011110100";
        wait for Clk_period; 
        Features_din <= "1111111010000001";
        wait for Clk_period; 
        Features_din <= "1111000110011011";
        wait for Clk_period; 
        Features_din <= "1111000011110111";
        wait for Clk_period; 
        Features_din <= "1111101010101011";
        wait for Clk_period; 
        Features_din <= "1111110100100001";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "1111011110110001";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001100000110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000000101100000";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "1111110110001000";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "0000001010011011";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011110101111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001001110000";
        wait for Clk_period; 
        Features_din <= "0000110101111000";
        wait for Clk_period; 
        Features_din <= "1111111000110101";
        wait for Clk_period; 
        Features_din <= "1111101111000011";
        wait for Clk_period; 
        Features_din <= "0000000011001101";
        wait for Clk_period; 
        Features_din <= "1111101100010001";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000100101101";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "1111111001001000";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000011001000011";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "1111111000010111";
        wait for Clk_period; 
        Features_din <= "1111100100111111";
        wait for Clk_period; 
        Features_din <= "0000001000011111";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "0000000110011110";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001000010010001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001001001011001";
        wait for Clk_period; 
        Features_din <= "0000010100100110";
        wait for Clk_period; 
        Features_din <= "1111011001100000";
        wait for Clk_period; 
        Features_din <= "1111110010001010";
        wait for Clk_period; 
        Features_din <= "1111110010100110";
        wait for Clk_period; 
        Features_din <= "1111010011101101";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000001001001011";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "1111110001000001";
        wait for Clk_period; 
        Features_din <= "1111100001011010";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000000111011010";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "0000010010100000";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000000110011100";
        wait for Clk_period; 
        Features_din <= "1111111111011000";
        wait for Clk_period; 
        Features_din <= "0000001000011000";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000001000110101";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000010111101";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000100100101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "1111110101000101";
        wait for Clk_period; 
        Features_din <= "0000101110010101";
        wait for Clk_period; 
        Features_din <= "0000001000101011";
        wait for Clk_period; 
        Features_din <= "1111110110010111";
        wait for Clk_period; 
        Features_din <= "1111010011111110";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "1111100111001100";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "0000001000101101";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111100111111010";
        wait for Clk_period; 
        Features_din <= "0000001100010011";
        wait for Clk_period; 
        Features_din <= "0000001010011010";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000011001010";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110000111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001010001011100";
        wait for Clk_period; 
        Features_din <= "0000001000000110";
        wait for Clk_period; 
        Features_din <= "1111011110001111";
        wait for Clk_period; 
        Features_din <= "1111111000100000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111010111011101";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000001011001000";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "1111110101000011";
        wait for Clk_period; 
        Features_din <= "1111101000110010";
        wait for Clk_period; 
        Features_din <= "0000001010001010";
        wait for Clk_period; 
        Features_din <= "0000001001111011";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "1111101110001101";
        wait for Clk_period; 
        Features_din <= "0000010011111101";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000000011101000";
        wait for Clk_period; 
        Features_din <= "0000000100111101";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000001011110101";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000011101001";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001111111111000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111101110101111";
        wait for Clk_period; 
        Features_din <= "1111111011000111";
        wait for Clk_period; 
        Features_din <= "1111100001111111";
        wait for Clk_period; 
        Features_din <= "1111100011101110";
        wait for Clk_period; 
        Features_din <= "0000010111111110";
        wait for Clk_period; 
        Features_din <= "1111010100110111";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "1111101010110110";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000000110110111";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "1111100110100111";
        wait for Clk_period; 
        Features_din <= "0000001001101010";
        wait for Clk_period; 
        Features_din <= "0000000110010111";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "0000000011000111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001110011010110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011011011";
        wait for Clk_period; 
        Features_din <= "1111111010011111";
        wait for Clk_period; 
        Features_din <= "1111001100001011";
        wait for Clk_period; 
        Features_din <= "1111010011110101";
        wait for Clk_period; 
        Features_din <= "1111101101000000";
        wait for Clk_period; 
        Features_din <= "1111101010000110";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000001011011010";
        wait for Clk_period; 
        Features_din <= "0000010010000001";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111110101111111";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000010100000010";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "1111111000100101";
        wait for Clk_period; 
        Features_din <= "1111100100011011";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000010111101";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001001000011000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010101111010";
        wait for Clk_period; 
        Features_din <= "0000000110100001";
        wait for Clk_period; 
        Features_din <= "1111011101111011";
        wait for Clk_period; 
        Features_din <= "1111110111010100";
        wait for Clk_period; 
        Features_din <= "1111101001110000";
        wait for Clk_period; 
        Features_din <= "1111011100001001";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "1111110010000000";
        wait for Clk_period; 
        Features_din <= "1111101011011010";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001011011100";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000000110100110";
        wait for Clk_period; 
        Features_din <= "1111101100110001";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000000101110100";
        wait for Clk_period; 
        Features_din <= "0000001010101100";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001110100011110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111111110100";
        wait for Clk_period; 
        Features_din <= "1111111101110110";
        wait for Clk_period; 
        Features_din <= "1111100101110001";
        wait for Clk_period; 
        Features_din <= "1111001011110010";
        wait for Clk_period; 
        Features_din <= "0000000111101111";
        wait for Clk_period; 
        Features_din <= "1111001010000010";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000001001010110";
        wait for Clk_period; 
        Features_din <= "0000010001110001";
        wait for Clk_period; 
        Features_din <= "0000001011110001";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000111001101";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "1111111001011010";
        wait for Clk_period; 
        Features_din <= "1111110110010101";
        wait for Clk_period; 
        Features_din <= "1111100001011100";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000001000000111";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "0000000010110011";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010101001001101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "1111001000101001";
        wait for Clk_period; 
        Features_din <= "1111001110001001";
        wait for Clk_period; 
        Features_din <= "1111101000011101";
        wait for Clk_period; 
        Features_din <= "1111000110110110";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111101001011111";
        wait for Clk_period; 
        Features_din <= "1111100110111011";
        wait for Clk_period; 
        Features_din <= "0000000110100100";
        wait for Clk_period; 
        Features_din <= "0000000111100111";
        wait for Clk_period; 
        Features_din <= "0000001011001110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010011000100";
        wait for Clk_period; 
        Features_din <= "0000001010010000";
        wait for Clk_period; 
        Features_din <= "0000000111110110";
        wait for Clk_period; 
        Features_din <= "1111111111001110";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000000011100100";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001010110010111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010001111101";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "1111101010010100";
        wait for Clk_period; 
        Features_din <= "1111010111011100";
        wait for Clk_period; 
        Features_din <= "1111110001010011";
        wait for Clk_period; 
        Features_din <= "1111100000111001";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000001011101011";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000000111110000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "1111111100011000";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "1111111010000101";
        wait for Clk_period; 
        Features_din <= "1111011110111000";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000000110001101";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001010111001011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010111011110";
        wait for Clk_period; 
        Features_din <= "0000011011111100";
        wait for Clk_period; 
        Features_din <= "1111100011001001";
        wait for Clk_period; 
        Features_din <= "1111101010111000";
        wait for Clk_period; 
        Features_din <= "1111110100100000";
        wait for Clk_period; 
        Features_din <= "1111010000110100";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000001100101000";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000001011011000";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000000110010011";
        wait for Clk_period; 
        Features_din <= "0000000111011001";
        wait for Clk_period; 
        Features_din <= "0000000101000011";
        wait for Clk_period; 
        Features_din <= "1111011011001010";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "0000000101001011";
        wait for Clk_period; 
        Features_din <= "1111111100000010";
        wait for Clk_period; 
        Features_din <= "0000000111100100";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001000000000101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000111000111001";
        wait for Clk_period; 
        Features_din <= "0000011011010110";
        wait for Clk_period; 
        Features_din <= "1111101000111101";
        wait for Clk_period; 
        Features_din <= "1111100101110001";
        wait for Clk_period; 
        Features_din <= "1111100101101110";
        wait for Clk_period; 
        Features_din <= "1111010011111101";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111101011101101";
        wait for Clk_period; 
        Features_din <= "0000010010110011";
        wait for Clk_period; 
        Features_din <= "0000000011111000";
        wait for Clk_period; 
        Features_din <= "0000001011001111";
        wait for Clk_period; 
        Features_din <= "0000001011000110";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111100101100101";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000000101101101";
        wait for Clk_period; 
        Features_din <= "1111111110000101";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001010111010";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000011010001";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001001100000111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000000101111000";
        wait for Clk_period; 
        Features_din <= "1111011101101101";
        wait for Clk_period; 
        Features_din <= "1111101111110001";
        wait for Clk_period; 
        Features_din <= "1111110000101111";
        wait for Clk_period; 
        Features_din <= "1111011010011111";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111101100000100";
        wait for Clk_period; 
        Features_din <= "1111100101011100";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000001000101000";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "0000010100001001";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000000110010110";
        wait for Clk_period; 
        Features_din <= "1111111110011111";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000011001110";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001101100000010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "1111001111011011";
        wait for Clk_period; 
        Features_din <= "1111011101000110";
        wait for Clk_period; 
        Features_din <= "1111101000101101";
        wait for Clk_period; 
        Features_din <= "1111101101101111";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111110011101000";
        wait for Clk_period; 
        Features_din <= "1111101011001101";
        wait for Clk_period; 
        Features_din <= "0000001000101111";
        wait for Clk_period; 
        Features_din <= "0000001100101001";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001001110001";
        wait for Clk_period; 
        Features_din <= "1111101011111111";
        wait for Clk_period; 
        Features_din <= "0000010011011001";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000000101100101";
        wait for Clk_period; 
        Features_din <= "0000001001110100";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000001001001100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001000000111010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "0001000100111001";
        wait for Clk_period; 
        Features_din <= "1111010011111010";
        wait for Clk_period; 
        Features_din <= "1111011100001110";
        wait for Clk_period; 
        Features_din <= "1111110111111000";
        wait for Clk_period; 
        Features_din <= "1111011010001110";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111101100001001";
        wait for Clk_period; 
        Features_din <= "1111100100111011";
        wait for Clk_period; 
        Features_din <= "0000001010110100";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000001010101100";
        wait for Clk_period; 
        Features_din <= "0000000110010000";
        wait for Clk_period; 
        Features_din <= "0000010011000111";
        wait for Clk_period; 
        Features_din <= "0000001011101111";
        wait for Clk_period; 
        Features_din <= "0000000110101110";
        wait for Clk_period; 
        Features_din <= "1111111110101011";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010010100001000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011001011101";
        wait for Clk_period; 
        Features_din <= "1111110111101011";
        wait for Clk_period; 
        Features_din <= "1110111000101100";
        wait for Clk_period; 
        Features_din <= "1111010110010001";
        wait for Clk_period; 
        Features_din <= "1111111001110010";
        wait for Clk_period; 
        Features_din <= "1111011011010100";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111101010001101";
        wait for Clk_period; 
        Features_din <= "1111100111001110";
        wait for Clk_period; 
        Features_din <= "0000001010010000";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001011010000";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000000100011001";
        wait for Clk_period; 
        Features_din <= "1111111101010101";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "0000000100111011";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010011101010001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000100100001110";
        wait for Clk_period; 
        Features_din <= "1111101101011100";
        wait for Clk_period; 
        Features_din <= "1110111111110010";
        wait for Clk_period; 
        Features_din <= "1111011111100110";
        wait for Clk_period; 
        Features_din <= "0000000101000110";
        wait for Clk_period; 
        Features_din <= "1111101101000111";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000011011001110";
        wait for Clk_period; 
        Features_din <= "1111110010001100";
        wait for Clk_period; 
        Features_din <= "0000000101001100";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "1111100111110101";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "1111110111010010";
        wait for Clk_period; 
        Features_din <= "0000000101001000";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "0000000011001110";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000110010011011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001010110011";
        wait for Clk_period; 
        Features_din <= "0000100011000110";
        wait for Clk_period; 
        Features_din <= "1111110011001101";
        wait for Clk_period; 
        Features_din <= "1111110010101000";
        wait for Clk_period; 
        Features_din <= "1111111111011101";
        wait for Clk_period; 
        Features_din <= "1111100100110010";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000011101011";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000100111001";
        wait for Clk_period; 
        Features_din <= "0000010011000010";
        wait for Clk_period; 
        Features_din <= "0000000111101110";
        wait for Clk_period; 
        Features_din <= "0000000101010000";
        wait for Clk_period; 
        Features_din <= "1111111000101000";
        wait for Clk_period; 
        Features_din <= "0000001010000001";
        wait for Clk_period; 
        Features_din <= "0000010110000111";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "1111111001101010";
        wait for Clk_period; 
        Features_din <= "1111100011100110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000001001110100";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "0000000011010010";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001111100010111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000101111000010";
        wait for Clk_period; 
        Features_din <= "0000101010100001";
        wait for Clk_period; 
        Features_din <= "1111000010011001";
        wait for Clk_period; 
        Features_din <= "1111011001001010";
        wait for Clk_period; 
        Features_din <= "1111101110000110";
        wait for Clk_period; 
        Features_din <= "1110100101110111";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000100100011";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000001010001000";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000100100011";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111011100101111";
        wait for Clk_period; 
        Features_din <= "0000000110101000";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "1111111000110100";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010001010111011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111110100011100";
        wait for Clk_period; 
        Features_din <= "0000001000011001";
        wait for Clk_period; 
        Features_din <= "1111010001100111";
        wait for Clk_period; 
        Features_din <= "1111000101010110";
        wait for Clk_period; 
        Features_din <= "1111110100101011";
        wait for Clk_period; 
        Features_din <= "1111011101001101";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000011111000";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000111110100";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000000100001110";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "1111100110000100";
        wait for Clk_period; 
        Features_din <= "0000001011110001";
        wait for Clk_period; 
        Features_din <= "1111101110100001";
        wait for Clk_period; 
        Features_din <= "1111110111001110";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000011001010";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001010010101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000000110011010";
        wait for Clk_period; 
        Features_din <= "0000010101100101";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "0000100011001011";
        wait for Clk_period; 
        Features_din <= "1111111011001001";
        wait for Clk_period; 
        Features_din <= "1111010110101101";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111011111000101";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "0000000110010011";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000000011101000";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "1111110110010001";
        wait for Clk_period; 
        Features_din <= "0000000110110000";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "0000001011000011";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "0000000011010001";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(3, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011000110111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001110010000100";
        wait for Clk_period; 
        Features_din <= "0000011101010111";
        wait for Clk_period; 
        Features_din <= "1111100011000010";
        wait for Clk_period; 
        Features_din <= "1111111001010010";
        wait for Clk_period; 
        Features_din <= "1111100011101000";
        wait for Clk_period; 
        Features_din <= "1110111000111100";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "1111100100110011";
        wait for Clk_period; 
        Features_din <= "1111111100010000";
        wait for Clk_period; 
        Features_din <= "0000000101110101";
        wait for Clk_period; 
        Features_din <= "0000000011010011";
        wait for Clk_period; 
        Features_din <= "0000011110111010";
        wait for Clk_period; 
        Features_din <= "0000000100111000";
        wait for Clk_period; 
        Features_din <= "0000000110010000";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "1111111011110110";
        wait for Clk_period; 
        Features_din <= "1111111011011110";
        wait for Clk_period; 
        Features_din <= "0000000100011000";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001000000101";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "0000000100100001";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(2, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011011111011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010010010100";
        wait for Clk_period; 
        Features_din <= "1111111000111110";
        wait for Clk_period; 
        Features_din <= "0000000100111010";
        wait for Clk_period; 
        Features_din <= "1111110011110110";
        wait for Clk_period; 
        Features_din <= "1111111010001010";
        wait for Clk_period; 
        Features_din <= "1111010011100101";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000110010010";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111110000001100";
        wait for Clk_period; 
        Features_din <= "1111101101000101";
        wait for Clk_period; 
        Features_din <= "0000000111011100";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000000101100000";
        wait for Clk_period; 
        Features_din <= "1111101100101010";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000000101111110";
        wait for Clk_period; 
        Features_din <= "0000000110010110";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001000101001";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000011111110";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010001101010100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011010110010";
        wait for Clk_period; 
        Features_din <= "1111111001110010";
        wait for Clk_period; 
        Features_din <= "1110111010000110";
        wait for Clk_period; 
        Features_din <= "1111101000111100";
        wait for Clk_period; 
        Features_din <= "1111101100010111";
        wait for Clk_period; 
        Features_din <= "1111000111110011";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000001000000001";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000010100011010";
        wait for Clk_period; 
        Features_din <= "1111101000010111";
        wait for Clk_period; 
        Features_din <= "0000001000111000";
        wait for Clk_period; 
        Features_din <= "0000000110010110";
        wait for Clk_period; 
        Features_din <= "1111111010101101";
        wait for Clk_period; 
        Features_din <= "0000000101010101";
        wait for Clk_period; 
        Features_din <= "0000010110110110";
        wait for Clk_period; 
        Features_din <= "1111110100111110";
        wait for Clk_period; 
        Features_din <= "1111110101111111";
        wait for Clk_period; 
        Features_din <= "0000000110101110";
        wait for Clk_period; 
        Features_din <= "0000001100010100";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000001100001101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000010111111";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001111011100111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000110101101000";
        wait for Clk_period; 
        Features_din <= "1111110000101101";
        wait for Clk_period; 
        Features_din <= "1111011000000100";
        wait for Clk_period; 
        Features_din <= "1111010111011101";
        wait for Clk_period; 
        Features_din <= "1111100101111110";
        wait for Clk_period; 
        Features_din <= "1111000111111110";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000011101111110";
        wait for Clk_period; 
        Features_din <= "1111101100000010";
        wait for Clk_period; 
        Features_din <= "0000000101101111";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "1111110000111001";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111111011010110";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000000110101110";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "0000000011010111";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001011101010111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111110101101110";
        wait for Clk_period; 
        Features_din <= "1111110011000011";
        wait for Clk_period; 
        Features_din <= "1111100010011001";
        wait for Clk_period; 
        Features_din <= "1111101011111101";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111100111101000";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "1111101100101011";
        wait for Clk_period; 
        Features_din <= "1111100100111111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000000111010110";
        wait for Clk_period; 
        Features_din <= "0000000110000000";
        wait for Clk_period; 
        Features_din <= "0000010100111101";
        wait for Clk_period; 
        Features_din <= "0000001011011010";
        wait for Clk_period; 
        Features_din <= "0000001000000000";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "0000000111001101";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "0000000011000101";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000011001111";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001101001010000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000100101011011";
        wait for Clk_period; 
        Features_din <= "1111111101100000";
        wait for Clk_period; 
        Features_din <= "1110111100010000";
        wait for Clk_period; 
        Features_din <= "1110111000100000";
        wait for Clk_period; 
        Features_din <= "1111110011100001";
        wait for Clk_period; 
        Features_din <= "1111010111010110";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000110010010";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111011101010111";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000000110101000";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000001011010100";
        wait for Clk_period; 
        Features_din <= "0000000100000110";
        wait for Clk_period; 
        Features_din <= "0000001011000111";
        wait for Clk_period; 
        Features_din <= "0000000110011001";
        wait for Clk_period; 
        Features_din <= "1111111110111001";
        wait for Clk_period; 
        Features_din <= "1111110111110000";
        wait for Clk_period; 
        Features_din <= "0000000110001101";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000000100000010";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "0000000010111110";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010010000111000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111110111000101";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "1110111001100001";
        wait for Clk_period; 
        Features_din <= "1111001101101100";
        wait for Clk_period; 
        Features_din <= "1111011101001000";
        wait for Clk_period; 
        Features_din <= "1111100001011010";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111110110000101";
        wait for Clk_period; 
        Features_din <= "1111111000001000";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000100110000000";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "1111110110000000";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "1111111000001000";
        wait for Clk_period; 
        Features_din <= "1111111011011100";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010001001000000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111101101110011";
        wait for Clk_period; 
        Features_din <= "1111111110011110";
        wait for Clk_period; 
        Features_din <= "1111001100101111";
        wait for Clk_period; 
        Features_din <= "1111101000111101";
        wait for Clk_period; 
        Features_din <= "1111110110011001";
        wait for Clk_period; 
        Features_din <= "1111011001000010";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "1111100111000111";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001100000100";
        wait for Clk_period; 
        Features_din <= "0000001010100011";
        wait for Clk_period; 
        Features_din <= "0000000111010101";
        wait for Clk_period; 
        Features_din <= "1111101000011100";
        wait for Clk_period; 
        Features_din <= "0000001100010000";
        wait for Clk_period; 
        Features_din <= "0000001000111011";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000001010100000";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "0000000010111000";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001111000111110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111011110011100";
        wait for Clk_period; 
        Features_din <= "1111011011111100";
        wait for Clk_period; 
        Features_din <= "1111100110110111";
        wait for Clk_period; 
        Features_din <= "1111100100100011";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111101100100101";
        wait for Clk_period; 
        Features_din <= "1111100110100011";
        wait for Clk_period; 
        Features_din <= "0000001010110100";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000000111001001";
        wait for Clk_period; 
        Features_din <= "0000000011011100";
        wait for Clk_period; 
        Features_din <= "0000011000010001";
        wait for Clk_period; 
        Features_din <= "0000001000111011";
        wait for Clk_period; 
        Features_din <= "0000000110100110";
        wait for Clk_period; 
        Features_din <= "1111111101111100";
        wait for Clk_period; 
        Features_din <= "0000001100010000";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000001011010010";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
            wait;
    end process;
end;
