

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.types.all;

entity image_test is
    generic(TREE_RAM_BITS: positive := 13;
            NUM_CLASSES:   positive := 8;
            NUM_FEATURES:  positive := 36);
end image_test;

architecture behavior of image_test is
    
    component image
        generic(TREE_RAM_BITS: positive;
                NUM_CLASSES:   positive;
                NUM_FEATURES:  positive);
        port(-- Control signals
             Clk:   in std_logic;
             Reset: in std_logic;
             
             -- Inputs for the nodes reception (trees)
             Load_trees: in std_logic;
             Valid_node: in std_logic;
             Addr:       in std_logic_vector(TREE_RAM_BITS - 1  downto 0);
             Trees_din:  in std_logic_vector(31 downto 0);
             
             -- Inputs for the features reception (pixels)
             Load_features: in std_logic;
             Valid_feature: in std_logic;
             Features_din:  in std_logic_vector(15 downto 0);
             Last_feature:  in std_logic;
             
             -- Output signals
             --     Finish:     finish (also 'ready') signal
             --     Dout:       the selected class
             --     Greater:    the value of the selected class prediction
             --     Curr_state: the current state
             Finish:     out std_logic;
             Dout:       out std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);
             greater:    out std_logic_vector(31 downto 0);
             curr_state: out std_logic_vector(2 downto 0));
    end component;
    
    component counter is
        generic(BITS: natural);
        port(Clk:   in  std_logic;
             Reset: in  std_logic;
             Count: in  std_logic;
             Dout:  out std_logic_vector (BITS - 1 downto 0));
    end component;
    
    -- Inputs
    signal Clk:           std_logic := '0';
    signal Reset:         std_logic := '0';
    signal Load_trees:    std_logic := '0';
    signal Valid_node:    std_logic := '0';
    signal Addr:          std_logic_vector(TREE_RAM_BITS - 1 downto
                                           0) := (others => '0');
    signal Trees_din:     std_logic_vector(31 downto 0) := (others => '0');
    signal Load_features: std_logic := '0';
    signal Valid_feature: std_logic := '0';
    signal Features_din:  std_logic_vector(15 downto 0) := (others => '0');
    signal last_feature:  std_logic := '0';
    
    -- Outputs
    signal Finish:     std_logic;
    signal Dout:       std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);
    signal greater:    std_logic_vector(31 downto 0);
    signal curr_state: std_logic_vector(2 downto 0);
    
    -- Clock period definition
    constant Clk_period : time := 10 ns;
    
    -- Counter signals
    signal pc_count, hc_count: std_logic := '0';
    signal pixels, hits: std_logic_vector(15 downto 0) := (others => '0');
    
    -- Label signal
    signal class_label: std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);

begin
    
    -- Instantiate the Unit Under Test (UUT)
    uut: image
        generic map(TREE_RAM_BITS => TREE_RAM_BITS,
                    NUM_CLASSES   => NUM_CLASSES,
                    NUM_FEATURES  => NUM_FEATURES)
        port map(Clk           => Clk,
                 Reset         => Reset,
                 Load_trees    => Load_trees,
                 Valid_node    => Valid_node,
                 Addr          => Addr,
                 Trees_din     => Trees_din,
                 Load_features => Load_features,
                 Valid_feature => Valid_feature,
                 Features_din  => Features_din,
                 Last_feature  => Last_feature,
                 Finish        => Finish,
                 Dout          => Dout,
                 greater       => greater,
                 curr_state    => curr_state);
    
    -- To count the pixels
    pixel_counter: counter
        generic map(BITS => 16)
        port map(Clk   => Clk, 
                 Reset => Reset,
                 Count => pc_count,
                 Dout  => pixels);
    
    -- To count the hits
    hit_counter: counter
        generic map(BITS => 16)
        port map(Clk   => Clk, 
                 Reset => Reset,
                 Count => hc_count,
                 Dout  => hits);
    
    -- Clock process definition
    Clk_process: process
    begin
        Clk <= '0';
        wait for Clk_period/2;
        Clk <= '1';
        wait for Clk_period/2;
    end process;
    
    -- Stimulus process
    stim_proc: process
    begin
        
        Reset <= '1';
        
        -- hold reset state for 100 ns.
        wait for 100 ns;
        
        Reset <= '0';
        
        wait for Clk_period*10;
        


        
        -- LOAD TREES
        -----------------------------------------------------------------------
        
        -- Load and valid trees flags
        Load_trees <= '1';
        Valid_node <= '1';

        -- Class  0
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"010b835c";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"010a0130";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"01063114";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"01039604";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"ff560185";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"05f98208";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"0d000504";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"00040185";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"ff640185";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"10004904";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"008d0185";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"ff610185";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"00090f10";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"05fb0008";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"06fc7d04";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"ffc20185";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"006e0185";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"06ff2a04";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"00000185";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"021b0185";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"1dfd4704";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"012b0185";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"05f9b704";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"ff820185";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"007f0185";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"000c8b1c";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"06fbd20c";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"0900e008";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"1302f104";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"ff8c0185";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"017d0185";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"ff7e0185";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"0b009408";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"09010404";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"02020185";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"ff9c0185";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"0004eb04";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"015c0185";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"ff790185";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"09005204";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"015c0185";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"0f000004";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"005b0185";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"000cf204";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"00210185";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"ff590185";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"000f1c34";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"010e5020";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"000b3310";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"070a0708";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"030a3b04";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"03780185";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"00700185";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"02ffd204";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"ff9c0185";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"00ca0185";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"17f76d08";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"0401b904";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"00440185";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"01ae0185";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"1afadd04";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"006c0185";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"025d0185";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"070b480c";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"01100908";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"000c7a04";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"04380185";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"023d0185";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"04970185";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"0d005804";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"022f0185";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"00210185";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"01107c20";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"010f8d10";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"06ff2a08";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"04fde904";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"00ca0185";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"ff650185";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"00126b04";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"00e10185";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"ff8b0185";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"04000308";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"06ff1504";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"ff7c0185";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"00df0185";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"00131c04";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"02370185";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"ff9c0185";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"00126b08";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"03f7c704";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"03f10185";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"01910185";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"01134408";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"0900c804";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"ff880185";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"00a90185";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"02eb0185";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"010a814c";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"01063120";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"01039604";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"ff5c02c9";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"05f98210";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"08003308";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"0c00bc04";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"ffb602c9";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"014302c9";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"13040004";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"ff6602c9";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"000f02c9";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"10004908";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"07ffd204";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"ffd802c9";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"00f802c9";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"ff6702c9";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"00090f1c";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"06fc7d0c";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"1b026b08";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"1afd4304";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"00a002c9";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"ff7202c9";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"ff6302c9";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"020ad308";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"0900ec04";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"008702c9";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"014f02c9";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"06046d04";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"ff6a02c9";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"006c02c9";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"1dfd4704";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"013202c9";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"00106808";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"03f47604";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"00da02c9";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"ffb702c9";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"ff5c02c9";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"000de228";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"010cb714";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"0a003a04";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"ff6502c9";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"06fb9c08";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"0900b304";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"017702c9";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"ffa702c9";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"0900e904";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"015e02c9";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"009f02c9";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"0111b010";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"0009cb08";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"14003404";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"000c02c9";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"01a202c9";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"0702a704";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"016502c9";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"ff9102c9";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"01b702c9";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"010f4120";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"0011a310";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"0e003108";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"0b006f04";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"ffd502c9";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"010802c9";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"010ed104";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"ff9302c9";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"00ed02c9";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"0d000108";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"00126b04";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"00ce02c9";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"ffa302c9";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"0601e804";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"ff5f02c9";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"002602c9";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"0017800c";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"01138808";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"00109804";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"016b02c9";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"008d02c9";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"01cc02c9";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"ff9002c9";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"010a0150";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"01052520";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"0103960c";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"04f80e08";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"08003b04";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"00460435";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"ff770435";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"ff5f0435";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"0900e308";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"19006504";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"ff5c0435";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"003e0435";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"06005d04";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"ff770435";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"06048d04";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"01880435";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"ff850435";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"00090f1c";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"0c00f110";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"06fd2508";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"01091704";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"ff860435";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"008b0435";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"04001f04";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"00690435";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"ffbf0435";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"05f7a708";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"05f48f04";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"003f0435";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"ff9a0435";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"01fa0435";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"1dfd4704";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"00a90435";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"05f91c08";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"06fbf104";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"009b0435";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"ff840435";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"04fdfc04";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"ff840435";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"014c0435";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"010ea63c";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"000d1b20";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"010b3c10";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"04fec108";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"04fcb604";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"009b0435";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"00060435";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"12008004";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"01390435";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"00250435";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"00099608";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"0a003c04";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"00650435";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"01190435";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"03faa404";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"00d10435";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"ffa50435";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"0011a310";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"06ff2008";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"08003e04";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"004f0435";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"ff6e0435";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"010c1204";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"ffb60435";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"01030435";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"0601f908";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"15003204";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"00140435";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"ff640435";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"001e0435";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"00131c18";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"0111c210";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"000f8608";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"0f03e804";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"011a0435";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"00230435";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"19000104";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"00eb0435";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"ffd80435";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"0b00b704";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"01360435";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"008c0435";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"0f001108";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"1403f804";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"002c0435";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"ff760435";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"00178008";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"0e002c04";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"016b0435";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"002d0435";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"ffa10435";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"010a0154";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"01041e1c";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"01032f0c";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"04f80e08";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"1b027d04";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"ff8605c1";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"004205c1";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"ff6105c1";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"0900ec0c";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"01035108";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"12007b04";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"ffa605c1";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"004605c1";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"ff6705c1";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"005005c1";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"00090f18";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"0307c210";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"0c00f108";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"04009f04";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"003905c1";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"ffa905c1";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"0f01b104";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"014805c1";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"ffa305c1";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"0a004d04";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"ff6705c1";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"000b05c1";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"0900d010";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"12006908";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"0a004604";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"ff8f05c1";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"00c205c1";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"10002e04";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"003e05c1";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"ff5e05c1";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"0d000b08";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"03f71204";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"ffbf05c1";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"010c05c1";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"0205b504";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"004c05c1";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"ff7b05c1";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"010ea63c";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"000d1b1c";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"1402f30c";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"0b005e04";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"ff6d05c1";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"1f052404";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"012305c1";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"ffda05c1";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"010b3c08";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"0f009904";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"007505c1";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"ff7a05c1";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"1af8c104";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"ff6605c1";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"00b305c1";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"06ff2010";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"08003e08";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"08003804";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"ffa105c1";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"008a05c1";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"1e020904";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"002505c1";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"ff6005c1";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"010c1208";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"09008104";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"00ab05c1";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"ff6305c1";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"02057e04";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"fff205c1";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"00f105c1";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"000c4218";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"0b00600c";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"01115a08";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"0b006004";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"00a905c1";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"ffa105c1";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"00f905c1";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"020a9c08";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"23000004";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"00f505c1";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"002105c1";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"003005c1";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"0111c210";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"03f6c208";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"06ff3f04";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"002905c1";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"00a505c1";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"07fcb204";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"00de05c1";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"ff6405c1";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"17f74e08";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"03f7a104";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"00be05c1";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"ffb905c1";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"02085304";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"00fd05c1";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"002e05c1";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"01091744";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"01041e20";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"01032f14";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"04f80e08";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"0f003d04";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"ff8e0735";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"00400735";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"17f71108";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"03f4de04";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"00470735";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"ff7b0735";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"ff600735";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"0900df04";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"ff6b0735";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"07fef104";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"ff880735";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"00dd0735";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"00106820";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"06ff6f10";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"0c00d608";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"1102c504";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"ff950735";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"00810735";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"1403f804";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"ffdd0735";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"01560735";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"0d000608";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"1afcee04";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"01370735";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"ffca0735";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"05f99f04";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"ffcf0735";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"006b0735";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"ff680735";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"010ea640";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"000f5420";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"010bc110";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"000c8b08";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"0a003b04";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"ff890735";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"006b0735";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"03f47604";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"00d70735";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"ff9c0735";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"0e003808";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"0e002204";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"00690735";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"00b40735";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"0206f804";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"007b0735";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"ffda0735";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"15003610";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"04001f08";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"0d011704";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"01920735";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"00240735";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"0d025c04";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"ffa90735";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"00c20735";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"14040008";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"0b005d04";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"003f0735";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"ff610735";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"0c00a704";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"ffbf0735";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"00f60735";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"000b571c";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"070b4810";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"0b006008";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"02077f04";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"00b20735";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"ffbb0735";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"23000004";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"00d30735";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"00150735";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"0e003f08";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"04f99b04";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"00f90735";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"ff9a0735";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"ff6f0735";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"0111250c";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"16009008";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"15004b04";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"00760735";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"ff460735";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"011a0735";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"14040008";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"0d017004";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"00d20735";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"00a20735";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"01134404";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"00220735";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"00d40735";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"01091738";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"01041e20";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"01032f14";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"04f80e08";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"0a003f04";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"003f0869";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"ff950869";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"17f71108";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"0c00b004";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"ff820869";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"00480869";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"ff620869";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"0900df04";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"ff6f0869";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"07fef104";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"ff8f0869";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"00b70869";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"00106814";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"0307c210";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"15005308";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"0a004304";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"002f0869";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"ffd40869";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"05f75104";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"01610869";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"002d0869";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"ff6e0869";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"ff6d0869";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"010eef28";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"00126b20";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"05f9b710";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"010b3c08";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"21000004";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"00410869";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"ff970869";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"05f14a04";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"ff7e0869";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"006c0869";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"06faeb08";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"08004204";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"00070869";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"ff9a0869";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"08002004";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"fff40869";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"00e00869";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"0601c204";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"ff6e0869";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"00450869";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"0111c220";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"000c7a10";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"0b006008";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"0e004004";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"ffc80869";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"008d0869";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"0f03d704";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"00af0869";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"00000869";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"1302b408";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"1b027a04";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"00810869";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"ff960869";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"0a005904";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"007c0869";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"ff6c0869";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"000e190c";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"0b00b708";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"0e001404";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"00430869";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"00c90869";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"002d0869";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"000e6808";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"05f24904";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"fef90869";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"008e0869";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"17f71a04";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"00200869";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"00ad0869";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"010b284c";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"01052520";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"0900e00c";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"020ce804";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"ff6209dd";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"04fead04";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"00d809dd";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"ff7709dd";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"01032f08";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"04f80e04";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"004209dd";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"ff6909dd";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"04fca304";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"ff7709dd";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"07fcbd04";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"ffad09dd";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"00f709dd";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"1600a720";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"000bff10";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"10005108";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"03f72004";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"008209dd";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"001b09dd";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"0700bc04";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"ffff09dd";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"ff5609dd";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"10004108";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"08003c04";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"ff9509dd";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"00a009dd";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"0d000004";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"008409dd";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"ff6b09dd";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"0a005004";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"fffd09dd";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"0000f704";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"002209dd";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"017009dd";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"01107c3c";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"0009961c";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"0b005e0c";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"0c009308";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"0d000604";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"ffe309dd";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"007609dd";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"ff3009dd";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"06003008";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"010d7004";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"004a09dd";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"008a09dd";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"0206cf04";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"00ca09dd";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"007709dd";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"1af94c10";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"0c00b408";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"000a2a04";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"007009dd";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"ff3c09dd";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"010bf004";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"ff9209dd";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"009909dd";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"07004508";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"02020604";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"ff9709dd";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"005509dd";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"1100b004";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"009609dd";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"ff5009dd";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"07f87a20";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"14040010";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"0f009408";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"0f000004";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"000109dd";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"00a709dd";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"06ffa804";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"ffe109dd";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"00b409dd";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"0a004808";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"0b005d04";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"005d09dd";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"ff6009dd";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"04007504";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"009d09dd";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"002909dd";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"0800500c";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"0b00b708";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"0111f804";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"009f09dd";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"00bb09dd";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"001409dd";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"0a005304";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"008809dd";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"ff9409dd";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"0107ec48";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"0103961c";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"04f80e08";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"10004004";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"00440b69";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"ff9d0b69";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"17f71108";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"10004404";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"00450b69";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"ff8e0b69";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"01032f04";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"ff660b69";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"15003504";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"00440b69";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"ff8c0b69";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"0900e51c";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"070b4810";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"13040008";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"10003604";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"00500b69";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"ff9a0b69";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"0600f304";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"ffc30b69";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"012c0b69";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"070d1308";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"11014304";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"00290b69";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"01590b69";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"ffa80b69";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"04067d0c";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"18001604";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"ff6a0b69";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"16006004";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"01010b69";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"00060b69";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"01230b69";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"010ea640";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"0a003c20";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"05f4f810";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"19000808";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"03f90f04";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"ff800b69";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"00b30b69";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"1f028404";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"00d20b69";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"00040b69";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"0203d108";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"15003c04";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"008e0b69";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"ffa10b69";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"0f013e04";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"ff080b69";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"ffe90b69";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"06ff1a10";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"07f79c08";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"0204af04";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"00850b69";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"ff740b69";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"04019a04";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"00220b69";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"009e0b69";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"0004c308";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"0604df04";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"00c10b69";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"ffdf0b69";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"ffff0b69";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"00580b69";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"0111c220";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"000c4210";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"0b006008";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"0e004004";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"ff980b69";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"00600b69";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"07047404";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"00900b69";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"004b0b69";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"16009008";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"03f73104";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"00140b69";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"00790b69";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"0206b904";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"00e80b69";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"00550b69";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"000e1910";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"08002408";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"08002204";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"008d0b69";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"ff7d0b69";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"070c0a04";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"00b00b69";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"001f0b69";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"000e6808";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"05f24904";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"ff1c0b69";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"00770b69";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"19000204";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"00590b69";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"00bc0b69";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"010bc148";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"01052520";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"0900e00c";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"020ce804";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"ff650ca9";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"04fe5404";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"00d70ca9";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"ff810ca9";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"01032f08";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"0900e104";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"002a0ca9";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"ff6e0ca9";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"19000108";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"19000004";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"fffb0ca9";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"01310ca9";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"ff7e0ca9";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"00106820";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"16009910";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"18000808";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"06078104";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"ff950ca9";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"00b70ca9";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"0f000104";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"007d0ca9";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"00100ca9";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"0d000908";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"04fb7f04";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"001a0ca9";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"01130ca9";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"010a5104";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"ff820ca9";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"00510ca9";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"09005f04";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"00330ca9";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"ff6e0ca9";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"0111c234";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"05f8bc20";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"0f000010";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"1afc0608";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"1403f804";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"002a0ca9";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"00c40ca9";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"21000004";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"00150ca9";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"ff3e0ca9";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"0900e908";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"1403ff04";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"004c0ca9";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"008b0ca9";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"1101af04";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"003e0ca9";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"ffae0ca9";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"00fdce08";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"0702a704";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"00930ca9";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"ff3e0ca9";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"0b005404";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"ffde0ca9";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"06f99c04";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"00110ca9";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"00ba0ca9";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"000e1910";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"08002408";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"08002204";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"00830ca9";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"ff850ca9";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"070c0a04";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"00a80ca9";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"001c0ca9";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"000e6808";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"05f24904";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"ff330ca9";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"006f0ca9";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"19000208";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"02035f04";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"00a20ca9";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"00140ca9";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"00b10ca9";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"010d0250";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"01041e1c";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"07039314";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"17f71108";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"03f62904";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"00480e15";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"ff980e15";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"01032f04";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"ff690e15";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"03fc1e04";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"ff7e0e15";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"00440e15";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"07047404";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"00630e15";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"ff8a0e15";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"0a003c18";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"05f46b0c";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"19000004";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"ff8b0e15";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"00082b04";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"00df0e15";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"00270e15";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"04fa3304";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"00520e15";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"1900bd04";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"ff4c0e15";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"00330e15";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"00106810";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"15003108";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"010c2404";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"00070e15";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"ff3a0e15";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"0c00e804";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"00230e15";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"00e70e15";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"1f024c08";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"1e024b04";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"ffd60e15";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"00ca0e15";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"ff6d0e15";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"0111c23c";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"16005d1c";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"18003f0c";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"05f1a604";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"ffa40e15";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"000f3604";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"00b80e15";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"01350e15";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"000fee08";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"010d5f04";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"00000e15";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"007d0e15";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"1101b804";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"ff690e15";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"00670e15";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"10004210";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"00090f08";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"0c00b104";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"ffe80e15";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"00aa0e15";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"02055504";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"ff310e15";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"fff00e15";
		wait for Clk_period;
		Addr <=  "0001101101001";
		Trees_din <= x"09005208";
		wait for Clk_period;
		Addr <=  "0001101101010";
		Trees_din <= x"19000004";
		wait for Clk_period;
		Addr <=  "0001101101011";
		Trees_din <= x"feed0e15";
		wait for Clk_period;
		Addr <=  "0001101101100";
		Trees_din <= x"00050e15";
		wait for Clk_period;
		Addr <=  "0001101101101";
		Trees_din <= x"0f000004";
		wait for Clk_period;
		Addr <=  "0001101101110";
		Trees_din <= x"00160e15";
		wait for Clk_period;
		Addr <=  "0001101101111";
		Trees_din <= x"00540e15";
		wait for Clk_period;
		Addr <=  "0001101110000";
		Trees_din <= x"000e1910";
		wait for Clk_period;
		Addr <=  "0001101110001";
		Trees_din <= x"08002408";
		wait for Clk_period;
		Addr <=  "0001101110010";
		Trees_din <= x"08002204";
		wait for Clk_period;
		Addr <=  "0001101110011";
		Trees_din <= x"00780e15";
		wait for Clk_period;
		Addr <=  "0001101110100";
		Trees_din <= x"ff8e0e15";
		wait for Clk_period;
		Addr <=  "0001101110101";
		Trees_din <= x"070c0a04";
		wait for Clk_period;
		Addr <=  "0001101110110";
		Trees_din <= x"00a20e15";
		wait for Clk_period;
		Addr <=  "0001101110111";
		Trees_din <= x"00180e15";
		wait for Clk_period;
		Addr <=  "0001101111000";
		Trees_din <= x"0b007010";
		wait for Clk_period;
		Addr <=  "0001101111001";
		Trees_din <= x"0b006808";
		wait for Clk_period;
		Addr <=  "0001101111010";
		Trees_din <= x"14040004";
		wait for Clk_period;
		Addr <=  "0001101111011";
		Trees_din <= x"009d0e15";
		wait for Clk_period;
		Addr <=  "0001101111100";
		Trees_din <= x"ffcc0e15";
		wait for Clk_period;
		Addr <=  "0001101111101";
		Trees_din <= x"04ff9104";
		wait for Clk_period;
		Addr <=  "0001101111110";
		Trees_din <= x"00200e15";
		wait for Clk_period;
		Addr <=  "0001101111111";
		Trees_din <= x"ff3a0e15";
		wait for Clk_period;
		Addr <=  "0001110000000";
		Trees_din <= x"17f71a04";
		wait for Clk_period;
		Addr <=  "0001110000001";
		Trees_din <= x"ff990e15";
		wait for Clk_period;
		Addr <=  "0001110000010";
		Trees_din <= x"05ef3e04";
		wait for Clk_period;
		Addr <=  "0001110000011";
		Trees_din <= x"00010e15";
		wait for Clk_period;
		Addr <=  "0001110000100";
		Trees_din <= x"009d0e15";
		wait for Clk_period;
		Addr <=  "0001110000101";
		Trees_din <= x"010eef54";
		wait for Clk_period;
		Addr <=  "0001110000110";
		Trees_din <= x"01063120";
		wait for Clk_period;
		Addr <=  "0001110000111";
		Trees_din <= x"10004918";
		wait for Clk_period;
		Addr <=  "0001110001000";
		Trees_din <= x"13040010";
		wait for Clk_period;
		Addr <=  "0001110001001";
		Trees_din <= x"07036e08";
		wait for Clk_period;
		Addr <=  "0001110001010";
		Trees_din <= x"0e002304";
		wait for Clk_period;
		Addr <=  "0001110001011";
		Trees_din <= x"00040f69";
		wait for Clk_period;
		Addr <=  "0001110001100";
		Trees_din <= x"ff8c0f69";
		wait for Clk_period;
		Addr <=  "0001110001101";
		Trees_din <= x"08003c04";
		wait for Clk_period;
		Addr <=  "0001110001110";
		Trees_din <= x"008b0f69";
		wait for Clk_period;
		Addr <=  "0001110001111";
		Trees_din <= x"ffb10f69";
		wait for Clk_period;
		Addr <=  "0001110010000";
		Trees_din <= x"0c00ac04";
		wait for Clk_period;
		Addr <=  "0001110010001";
		Trees_din <= x"00120f69";
		wait for Clk_period;
		Addr <=  "0001110010010";
		Trees_din <= x"01080f69";
		wait for Clk_period;
		Addr <=  "0001110010011";
		Trees_din <= x"09012704";
		wait for Clk_period;
		Addr <=  "0001110010100";
		Trees_din <= x"ff660f69";
		wait for Clk_period;
		Addr <=  "0001110010101";
		Trees_din <= x"002a0f69";
		wait for Clk_period;
		Addr <=  "0001110010110";
		Trees_din <= x"14022714";
		wait for Clk_period;
		Addr <=  "0001110010111";
		Trees_din <= x"08002b08";
		wait for Clk_period;
		Addr <=  "0001110011000";
		Trees_din <= x"00068c04";
		wait for Clk_period;
		Addr <=  "0001110011001";
		Trees_din <= x"00100f69";
		wait for Clk_period;
		Addr <=  "0001110011010";
		Trees_din <= x"ff6b0f69";
		wait for Clk_period;
		Addr <=  "0001110011011";
		Trees_din <= x"04030208";
		wait for Clk_period;
		Addr <=  "0001110011100";
		Trees_din <= x"16006f04";
		wait for Clk_period;
		Addr <=  "0001110011101";
		Trees_din <= x"00c20f69";
		wait for Clk_period;
		Addr <=  "0001110011110";
		Trees_din <= x"00420f69";
		wait for Clk_period;
		Addr <=  "0001110011111";
		Trees_din <= x"ff970f69";
		wait for Clk_period;
		Addr <=  "0001110100000";
		Trees_din <= x"1600a710";
		wait for Clk_period;
		Addr <=  "0001110100001";
		Trees_din <= x"21002508";
		wait for Clk_period;
		Addr <=  "0001110100010";
		Trees_din <= x"10005604";
		wait for Clk_period;
		Addr <=  "0001110100011";
		Trees_din <= x"001c0f69";
		wait for Clk_period;
		Addr <=  "0001110100100";
		Trees_din <= x"ffc40f69";
		wait for Clk_period;
		Addr <=  "0001110100101";
		Trees_din <= x"02068c04";
		wait for Clk_period;
		Addr <=  "0001110100110";
		Trees_din <= x"ff620f69";
		wait for Clk_period;
		Addr <=  "0001110100111";
		Trees_din <= x"000d0f69";
		wait for Clk_period;
		Addr <=  "0001110101000";
		Trees_din <= x"12004c08";
		wait for Clk_period;
		Addr <=  "0001110101001";
		Trees_din <= x"04fb1404";
		wait for Clk_period;
		Addr <=  "0001110101010";
		Trees_din <= x"008c0f69";
		wait for Clk_period;
		Addr <=  "0001110101011";
		Trees_din <= x"ff5e0f69";
		wait for Clk_period;
		Addr <=  "0001110101100";
		Trees_din <= x"04fc1204";
		wait for Clk_period;
		Addr <=  "0001110101101";
		Trees_din <= x"00190f69";
		wait for Clk_period;
		Addr <=  "0001110101110";
		Trees_din <= x"00e00f69";
		wait for Clk_period;
		Addr <=  "0001110101111";
		Trees_din <= x"0111c230";
		wait for Clk_period;
		Addr <=  "0001110110000";
		Trees_din <= x"00075718";
		wait for Clk_period;
		Addr <=  "0001110110001";
		Trees_din <= x"0702eb08";
		wait for Clk_period;
		Addr <=  "0001110110010";
		Trees_din <= x"12005a04";
		wait for Clk_period;
		Addr <=  "0001110110011";
		Trees_din <= x"ffe40f69";
		wait for Clk_period;
		Addr <=  "0001110110100";
		Trees_din <= x"00a70f69";
		wait for Clk_period;
		Addr <=  "0001110110101";
		Trees_din <= x"0900e008";
		wait for Clk_period;
		Addr <=  "0001110110110";
		Trees_din <= x"0707e004";
		wait for Clk_period;
		Addr <=  "0001110110111";
		Trees_din <= x"009b0f69";
		wait for Clk_period;
		Addr <=  "0001110111000";
		Trees_din <= x"00010f69";
		wait for Clk_period;
		Addr <=  "0001110111001";
		Trees_din <= x"11019d04";
		wait for Clk_period;
		Addr <=  "0001110111010";
		Trees_din <= x"00530f69";
		wait for Clk_period;
		Addr <=  "0001110111011";
		Trees_din <= x"ff0a0f69";
		wait for Clk_period;
		Addr <=  "0001110111100";
		Trees_din <= x"0a005a10";
		wait for Clk_period;
		Addr <=  "0001110111101";
		Trees_din <= x"0b006408";
		wait for Clk_period;
		Addr <=  "0001110111110";
		Trees_din <= x"0e003e04";
		wait for Clk_period;
		Addr <=  "0001110111111";
		Trees_din <= x"ff6b0f69";
		wait for Clk_period;
		Addr <=  "0001111000000";
		Trees_din <= x"00340f69";
		wait for Clk_period;
		Addr <=  "0001111000001";
		Trees_din <= x"03f77504";
		wait for Clk_period;
		Addr <=  "0001111000010";
		Trees_din <= x"00240f69";
		wait for Clk_period;
		Addr <=  "0001111000011";
		Trees_din <= x"00700f69";
		wait for Clk_period;
		Addr <=  "0001111000100";
		Trees_din <= x"16007404";
		wait for Clk_period;
		Addr <=  "0001111000101";
		Trees_din <= x"ff0c0f69";
		wait for Clk_period;
		Addr <=  "0001111000110";
		Trees_din <= x"001c0f69";
		wait for Clk_period;
		Addr <=  "0001111000111";
		Trees_din <= x"000e1914";
		wait for Clk_period;
		Addr <=  "0001111001000";
		Trees_din <= x"08002408";
		wait for Clk_period;
		Addr <=  "0001111001001";
		Trees_din <= x"08002204";
		wait for Clk_period;
		Addr <=  "0001111001010";
		Trees_din <= x"00700f69";
		wait for Clk_period;
		Addr <=  "0001111001011";
		Trees_din <= x"ff970f69";
		wait for Clk_period;
		Addr <=  "0001111001100";
		Trees_din <= x"070c0a08";
		wait for Clk_period;
		Addr <=  "0001111001101";
		Trees_din <= x"08003004";
		wait for Clk_period;
		Addr <=  "0001111001110";
		Trees_din <= x"005c0f69";
		wait for Clk_period;
		Addr <=  "0001111001111";
		Trees_din <= x"009f0f69";
		wait for Clk_period;
		Addr <=  "0001111010000";
		Trees_din <= x"00170f69";
		wait for Clk_period;
		Addr <=  "0001111010001";
		Trees_din <= x"000e6808";
		wait for Clk_period;
		Addr <=  "0001111010010";
		Trees_din <= x"05f24904";
		wait for Clk_period;
		Addr <=  "0001111010011";
		Trees_din <= x"ff490f69";
		wait for Clk_period;
		Addr <=  "0001111010100";
		Trees_din <= x"00630f69";
		wait for Clk_period;
		Addr <=  "0001111010101";
		Trees_din <= x"0900aa04";
		wait for Clk_period;
		Addr <=  "0001111010110";
		Trees_din <= x"00a10f69";
		wait for Clk_period;
		Addr <=  "0001111010111";
		Trees_din <= x"02035f04";
		wait for Clk_period;
		Addr <=  "0001111011000";
		Trees_din <= x"008e0f69";
		wait for Clk_period;
		Addr <=  "0001111011001";
		Trees_din <= x"fffe0f69";
		wait for Clk_period;
		Addr <=  "0001111011010";
		Trees_din <= x"010eef5c";
		wait for Clk_period;
		Addr <=  "0001111011011";
		Trees_din <= x"01054b24";
		wait for Clk_period;
		Addr <=  "0001111011100";
		Trees_din <= x"15003914";
		wait for Clk_period;
		Addr <=  "0001111011101";
		Trees_din <= x"18001c08";
		wait for Clk_period;
		Addr <=  "0001111011110";
		Trees_din <= x"03f78d04";
		wait for Clk_period;
		Addr <=  "0001111011111";
		Trees_din <= x"00ef10ed";
		wait for Clk_period;
		Addr <=  "0001111100000";
		Trees_din <= x"ffd710ed";
		wait for Clk_period;
		Addr <=  "0001111100001";
		Trees_din <= x"00036a08";
		wait for Clk_period;
		Addr <=  "0001111100010";
		Trees_din <= x"16005b04";
		wait for Clk_period;
		Addr <=  "0001111100011";
		Trees_din <= x"ffb410ed";
		wait for Clk_period;
		Addr <=  "0001111100100";
		Trees_din <= x"008b10ed";
		wait for Clk_period;
		Addr <=  "0001111100101";
		Trees_din <= x"ff7410ed";
		wait for Clk_period;
		Addr <=  "0001111100110";
		Trees_din <= x"0900e404";
		wait for Clk_period;
		Addr <=  "0001111100111";
		Trees_din <= x"ff6910ed";
		wait for Clk_period;
		Addr <=  "0001111101000";
		Trees_din <= x"0900e504";
		wait for Clk_period;
		Addr <=  "0001111101001";
		Trees_din <= x"008110ed";
		wait for Clk_period;
		Addr <=  "0001111101010";
		Trees_din <= x"0204af04";
		wait for Clk_period;
		Addr <=  "0001111101011";
		Trees_din <= x"ffef10ed";
		wait for Clk_period;
		Addr <=  "0001111101100";
		Trees_din <= x"ff7810ed";
		wait for Clk_period;
		Addr <=  "0001111101101";
		Trees_din <= x"14022718";
		wait for Clk_period;
		Addr <=  "0001111101110";
		Trees_din <= x"1dfd620c";
		wait for Clk_period;
		Addr <=  "0001111101111";
		Trees_din <= x"19000708";
		wait for Clk_period;
		Addr <=  "0001111110000";
		Trees_din <= x"07fd9f04";
		wait for Clk_period;
		Addr <=  "0001111110001";
		Trees_din <= x"ffeb10ed";
		wait for Clk_period;
		Addr <=  "0001111110010";
		Trees_din <= x"00b710ed";
		wait for Clk_period;
		Addr <=  "0001111110011";
		Trees_din <= x"011a10ed";
		wait for Clk_period;
		Addr <=  "0001111110100";
		Trees_din <= x"03f5d504";
		wait for Clk_period;
		Addr <=  "0001111110101";
		Trees_din <= x"ff7110ed";
		wait for Clk_period;
		Addr <=  "0001111110110";
		Trees_din <= x"010a1304";
		wait for Clk_period;
		Addr <=  "0001111110111";
		Trees_din <= x"ffcf10ed";
		wait for Clk_period;
		Addr <=  "0001111111000";
		Trees_din <= x"008310ed";
		wait for Clk_period;
		Addr <=  "0001111111001";
		Trees_din <= x"04020710";
		wait for Clk_period;
		Addr <=  "0001111111010";
		Trees_din <= x"07f7b808";
		wait for Clk_period;
		Addr <=  "0001111111011";
		Trees_din <= x"03f9bb04";
		wait for Clk_period;
		Addr <=  "0001111111100";
		Trees_din <= x"ffa010ed";
		wait for Clk_period;
		Addr <=  "0001111111101";
		Trees_din <= x"006810ed";
		wait for Clk_period;
		Addr <=  "0001111111110";
		Trees_din <= x"05f37304";
		wait for Clk_period;
		Addr <=  "0001111111111";
		Trees_din <= x"004e10ed";
		wait for Clk_period;
		Addr <=  "0010000000000";
		Trees_din <= x"000710ed";
		wait for Clk_period;
		Addr <=  "0010000000001";
		Trees_din <= x"0d008d08";
		wait for Clk_period;
		Addr <=  "0010000000010";
		Trees_din <= x"17f72e04";
		wait for Clk_period;
		Addr <=  "0010000000011";
		Trees_din <= x"ffe610ed";
		wait for Clk_period;
		Addr <=  "0010000000100";
		Trees_din <= x"009010ed";
		wait for Clk_period;
		Addr <=  "0010000000101";
		Trees_din <= x"010ab104";
		wait for Clk_period;
		Addr <=  "0010000000110";
		Trees_din <= x"ff7210ed";
		wait for Clk_period;
		Addr <=  "0010000000111";
		Trees_din <= x"002210ed";
		wait for Clk_period;
		Addr <=  "0010000001000";
		Trees_din <= x"0111c238";
		wait for Clk_period;
		Addr <=  "0010000001001";
		Trees_din <= x"00075718";
		wait for Clk_period;
		Addr <=  "0010000001010";
		Trees_din <= x"0702eb08";
		wait for Clk_period;
		Addr <=  "0010000001011";
		Trees_din <= x"12005a04";
		wait for Clk_period;
		Addr <=  "0010000001100";
		Trees_din <= x"ffdf10ed";
		wait for Clk_period;
		Addr <=  "0010000001101";
		Trees_din <= x"00a310ed";
		wait for Clk_period;
		Addr <=  "0010000001110";
		Trees_din <= x"04fa6808";
		wait for Clk_period;
		Addr <=  "0010000001111";
		Trees_din <= x"0e004504";
		wait for Clk_period;
		Addr <=  "0010000010000";
		Trees_din <= x"009510ed";
		wait for Clk_period;
		Addr <=  "0010000010001";
		Trees_din <= x"000210ed";
		wait for Clk_period;
		Addr <=  "0010000010010";
		Trees_din <= x"0c00b304";
		wait for Clk_period;
		Addr <=  "0010000010011";
		Trees_din <= x"ff8810ed";
		wait for Clk_period;
		Addr <=  "0010000010100";
		Trees_din <= x"008510ed";
		wait for Clk_period;
		Addr <=  "0010000010101";
		Trees_din <= x"04fd5410";
		wait for Clk_period;
		Addr <=  "0010000010110";
		Trees_din <= x"0e003b08";
		wait for Clk_period;
		Addr <=  "0010000010111";
		Trees_din <= x"0c00b904";
		wait for Clk_period;
		Addr <=  "0010000011000";
		Trees_din <= x"007410ed";
		wait for Clk_period;
		Addr <=  "0010000011001";
		Trees_din <= x"ffc210ed";
		wait for Clk_period;
		Addr <=  "0010000011010";
		Trees_din <= x"01108f04";
		wait for Clk_period;
		Addr <=  "0010000011011";
		Trees_din <= x"fefc10ed";
		wait for Clk_period;
		Addr <=  "0010000011100";
		Trees_din <= x"003410ed";
		wait for Clk_period;
		Addr <=  "0010000011101";
		Trees_din <= x"03f7ad08";
		wait for Clk_period;
		Addr <=  "0010000011110";
		Trees_din <= x"10004204";
		wait for Clk_period;
		Addr <=  "0010000011111";
		Trees_din <= x"ffda10ed";
		wait for Clk_period;
		Addr <=  "0010000100000";
		Trees_din <= x"004410ed";
		wait for Clk_period;
		Addr <=  "0010000100001";
		Trees_din <= x"17f7a404";
		wait for Clk_period;
		Addr <=  "0010000100010";
		Trees_din <= x"001510ed";
		wait for Clk_period;
		Addr <=  "0010000100011";
		Trees_din <= x"00a710ed";
		wait for Clk_period;
		Addr <=  "0010000100100";
		Trees_din <= x"000e1914";
		wait for Clk_period;
		Addr <=  "0010000100101";
		Trees_din <= x"08002408";
		wait for Clk_period;
		Addr <=  "0010000100110";
		Trees_din <= x"08002204";
		wait for Clk_period;
		Addr <=  "0010000100111";
		Trees_din <= x"006810ed";
		wait for Clk_period;
		Addr <=  "0010000101000";
		Trees_din <= x"ff9e10ed";
		wait for Clk_period;
		Addr <=  "0010000101001";
		Trees_din <= x"04f68e04";
		wait for Clk_period;
		Addr <=  "0010000101010";
		Trees_din <= x"002e10ed";
		wait for Clk_period;
		Addr <=  "0010000101011";
		Trees_din <= x"08003004";
		wait for Clk_period;
		Addr <=  "0010000101100";
		Trees_din <= x"005610ed";
		wait for Clk_period;
		Addr <=  "0010000101101";
		Trees_din <= x"009b10ed";
		wait for Clk_period;
		Addr <=  "0010000101110";
		Trees_din <= x"0b007010";
		wait for Clk_period;
		Addr <=  "0010000101111";
		Trees_din <= x"0b006808";
		wait for Clk_period;
		Addr <=  "0010000110000";
		Trees_din <= x"14040004";
		wait for Clk_period;
		Addr <=  "0010000110001";
		Trees_din <= x"008f10ed";
		wait for Clk_period;
		Addr <=  "0010000110010";
		Trees_din <= x"ffc610ed";
		wait for Clk_period;
		Addr <=  "0010000110011";
		Trees_din <= x"02044604";
		wait for Clk_period;
		Addr <=  "0010000110100";
		Trees_din <= x"003610ed";
		wait for Clk_period;
		Addr <=  "0010000110101";
		Trees_din <= x"ff5710ed";
		wait for Clk_period;
		Addr <=  "0010000110110";
		Trees_din <= x"17f71a04";
		wait for Clk_period;
		Addr <=  "0010000110111";
		Trees_din <= x"ffa210ed";
		wait for Clk_period;
		Addr <=  "0010000111000";
		Trees_din <= x"0600e104";
		wait for Clk_period;
		Addr <=  "0010000111001";
		Trees_din <= x"008e10ed";
		wait for Clk_period;
		Addr <=  "0010000111010";
		Trees_din <= x"fffb10ed";
		wait for Clk_period;
		Addr <=  "0010000111011";
		Trees_din <= x"0111b064";
		wait for Clk_period;
		Addr <=  "0010000111100";
		Trees_din <= x"0106bc24";
		wait for Clk_period;
		Addr <=  "0010000111101";
		Trees_din <= x"01032f0c";
		wait for Clk_period;
		Addr <=  "0010000111110";
		Trees_din <= x"04f80e04";
		wait for Clk_period;
		Addr <=  "0010000111111";
		Trees_din <= x"00261219";
		wait for Clk_period;
		Addr <=  "0010001000000";
		Trees_din <= x"17f71104";
		wait for Clk_period;
		Addr <=  "0010001000001";
		Trees_din <= x"000a1219";
		wait for Clk_period;
		Addr <=  "0010001000010";
		Trees_din <= x"ff6d1219";
		wait for Clk_period;
		Addr <=  "0010001000011";
		Trees_din <= x"020ce810";
		wait for Clk_period;
		Addr <=  "0010001000100";
		Trees_din <= x"0b007208";
		wait for Clk_period;
		Addr <=  "0010001000101";
		Trees_din <= x"0b006704";
		wait for Clk_period;
		Addr <=  "0010001000110";
		Trees_din <= x"ffe61219";
		wait for Clk_period;
		Addr <=  "0010001000111";
		Trees_din <= x"ff601219";
		wait for Clk_period;
		Addr <=  "0010001001000";
		Trees_din <= x"12007304";
		wait for Clk_period;
		Addr <=  "0010001001001";
		Trees_din <= x"00a41219";
		wait for Clk_period;
		Addr <=  "0010001001010";
		Trees_din <= x"ffe01219";
		wait for Clk_period;
		Addr <=  "0010001001011";
		Trees_din <= x"0900e404";
		wait for Clk_period;
		Addr <=  "0010001001100";
		Trees_din <= x"fffb1219";
		wait for Clk_period;
		Addr <=  "0010001001101";
		Trees_din <= x"011a1219";
		wait for Clk_period;
		Addr <=  "0010001001110";
		Trees_din <= x"0601ac20";
		wait for Clk_period;
		Addr <=  "0010001001111";
		Trees_din <= x"17f74210";
		wait for Clk_period;
		Addr <=  "0010001010000";
		Trees_din <= x"1b024608";
		wait for Clk_period;
		Addr <=  "0010001010001";
		Trees_din <= x"04ffbc04";
		wait for Clk_period;
		Addr <=  "0010001010010";
		Trees_din <= x"004e1219";
		wait for Clk_period;
		Addr <=  "0010001010011";
		Trees_din <= x"ffca1219";
		wait for Clk_period;
		Addr <=  "0010001010100";
		Trees_din <= x"03f6c204";
		wait for Clk_period;
		Addr <=  "0010001010101";
		Trees_din <= x"00281219";
		wait for Clk_period;
		Addr <=  "0010001010110";
		Trees_din <= x"ff9e1219";
		wait for Clk_period;
		Addr <=  "0010001010111";
		Trees_din <= x"16009108";
		wait for Clk_period;
		Addr <=  "0010001011000";
		Trees_din <= x"10005504";
		wait for Clk_period;
		Addr <=  "0010001011001";
		Trees_din <= x"001b1219";
		wait for Clk_period;
		Addr <=  "0010001011010";
		Trees_din <= x"ff871219";
		wait for Clk_period;
		Addr <=  "0010001011011";
		Trees_din <= x"0c007f04";
		wait for Clk_period;
		Addr <=  "0010001011100";
		Trees_din <= x"00921219";
		wait for Clk_period;
		Addr <=  "0010001011101";
		Trees_din <= x"00241219";
		wait for Clk_period;
		Addr <=  "0010001011110";
		Trees_din <= x"1c025c10";
		wait for Clk_period;
		Addr <=  "0010001011111";
		Trees_din <= x"10004608";
		wait for Clk_period;
		Addr <=  "0010001100000";
		Trees_din <= x"0c00a504";
		wait for Clk_period;
		Addr <=  "0010001100001";
		Trees_din <= x"ff671219";
		wait for Clk_period;
		Addr <=  "0010001100010";
		Trees_din <= x"005d1219";
		wait for Clk_period;
		Addr <=  "0010001100011";
		Trees_din <= x"08003604";
		wait for Clk_period;
		Addr <=  "0010001100100";
		Trees_din <= x"fffa1219";
		wait for Clk_period;
		Addr <=  "0010001100101";
		Trees_din <= x"00c11219";
		wait for Clk_period;
		Addr <=  "0010001100110";
		Trees_din <= x"05f7ca08";
		wait for Clk_period;
		Addr <=  "0010001100111";
		Trees_din <= x"010a0104";
		wait for Clk_period;
		Addr <=  "0010001101000";
		Trees_din <= x"ff8f1219";
		wait for Clk_period;
		Addr <=  "0010001101001";
		Trees_din <= x"002d1219";
		wait for Clk_period;
		Addr <=  "0010001101010";
		Trees_din <= x"0a003e04";
		wait for Clk_period;
		Addr <=  "0010001101011";
		Trees_din <= x"ffcd1219";
		wait for Clk_period;
		Addr <=  "0010001101100";
		Trees_din <= x"00b41219";
		wait for Clk_period;
		Addr <=  "0010001101101";
		Trees_din <= x"000e1918";
		wait for Clk_period;
		Addr <=  "0010001101110";
		Trees_din <= x"0b00a710";
		wait for Clk_period;
		Addr <=  "0010001101111";
		Trees_din <= x"04f68e04";
		wait for Clk_period;
		Addr <=  "0010001110000";
		Trees_din <= x"00281219";
		wait for Clk_period;
		Addr <=  "0010001110001";
		Trees_din <= x"000bb504";
		wait for Clk_period;
		Addr <=  "0010001110010";
		Trees_din <= x"009e1219";
		wait for Clk_period;
		Addr <=  "0010001110011";
		Trees_din <= x"03f7a104";
		wait for Clk_period;
		Addr <=  "0010001110100";
		Trees_din <= x"00941219";
		wait for Clk_period;
		Addr <=  "0010001110101";
		Trees_din <= x"ffd41219";
		wait for Clk_period;
		Addr <=  "0010001110110";
		Trees_din <= x"17f7fb04";
		wait for Clk_period;
		Addr <=  "0010001110111";
		Trees_din <= x"ff821219";
		wait for Clk_period;
		Addr <=  "0010001111000";
		Trees_din <= x"00681219";
		wait for Clk_period;
		Addr <=  "0010001111001";
		Trees_din <= x"0a004814";
		wait for Clk_period;
		Addr <=  "0010001111010";
		Trees_din <= x"0a004710";
		wait for Clk_period;
		Addr <=  "0010001111011";
		Trees_din <= x"1403fb08";
		wait for Clk_period;
		Addr <=  "0010001111100";
		Trees_din <= x"0f008d04";
		wait for Clk_period;
		Addr <=  "0010001111101";
		Trees_din <= x"009c1219";
		wait for Clk_period;
		Addr <=  "0010001111110";
		Trees_din <= x"fffa1219";
		wait for Clk_period;
		Addr <=  "0010001111111";
		Trees_din <= x"0203b504";
		wait for Clk_period;
		Addr <=  "0010010000000";
		Trees_din <= x"00611219";
		wait for Clk_period;
		Addr <=  "0010010000001";
		Trees_din <= x"ff701219";
		wait for Clk_period;
		Addr <=  "0010010000010";
		Trees_din <= x"ff5b1219";
		wait for Clk_period;
		Addr <=  "0010010000011";
		Trees_din <= x"12007004";
		wait for Clk_period;
		Addr <=  "0010010000100";
		Trees_din <= x"fffd1219";
		wait for Clk_period;
		Addr <=  "0010010000101";
		Trees_din <= x"00961219";
		wait for Clk_period;
		Addr <=  "0010010000110";
		Trees_din <= x"0111b04c";
		wait for Clk_period;
		Addr <=  "0010010000111";
		Trees_din <= x"01032f0c";
		wait for Clk_period;
		Addr <=  "0010010001000";
		Trees_din <= x"04f80e04";
		wait for Clk_period;
		Addr <=  "0010010001001";
		Trees_din <= x"0025131d";
		wait for Clk_period;
		Addr <=  "0010010001010";
		Trees_din <= x"17f71104";
		wait for Clk_period;
		Addr <=  "0010010001011";
		Trees_din <= x"000f131d";
		wait for Clk_period;
		Addr <=  "0010010001100";
		Trees_din <= x"ff70131d";
		wait for Clk_period;
		Addr <=  "0010010001101";
		Trees_din <= x"010bc120";
		wait for Clk_period;
		Addr <=  "0010010001110";
		Trees_din <= x"0f000110";
		wait for Clk_period;
		Addr <=  "0010010001111";
		Trees_din <= x"03f8cb08";
		wait for Clk_period;
		Addr <=  "0010010010000";
		Trees_din <= x"06fd6e04";
		wait for Clk_period;
		Addr <=  "0010010010001";
		Trees_din <= x"0160131d";
		wait for Clk_period;
		Addr <=  "0010010010010";
		Trees_din <= x"0045131d";
		wait for Clk_period;
		Addr <=  "0010010010011";
		Trees_din <= x"0b007604";
		wait for Clk_period;
		Addr <=  "0010010010100";
		Trees_din <= x"0033131d";
		wait for Clk_period;
		Addr <=  "0010010010101";
		Trees_din <= x"ff80131d";
		wait for Clk_period;
		Addr <=  "0010010010110";
		Trees_din <= x"0c00e608";
		wait for Clk_period;
		Addr <=  "0010010010111";
		Trees_din <= x"0a003d04";
		wait for Clk_period;
		Addr <=  "0010010011000";
		Trees_din <= x"ff9c131d";
		wait for Clk_period;
		Addr <=  "0010010011001";
		Trees_din <= x"fff8131d";
		wait for Clk_period;
		Addr <=  "0010010011010";
		Trees_din <= x"05f7fb04";
		wait for Clk_period;
		Addr <=  "0010010011011";
		Trees_din <= x"000f131d";
		wait for Clk_period;
		Addr <=  "0010010011100";
		Trees_din <= x"00ad131d";
		wait for Clk_period;
		Addr <=  "0010010011101";
		Trees_din <= x"05f8bc10";
		wait for Clk_period;
		Addr <=  "0010010011110";
		Trees_din <= x"0e003808";
		wait for Clk_period;
		Addr <=  "0010010011111";
		Trees_din <= x"0900e904";
		wait for Clk_period;
		Addr <=  "0010010100000";
		Trees_din <= x"0031131d";
		wait for Clk_period;
		Addr <=  "0010010100001";
		Trees_din <= x"fffd131d";
		wait for Clk_period;
		Addr <=  "0010010100010";
		Trees_din <= x"04fee704";
		wait for Clk_period;
		Addr <=  "0010010100011";
		Trees_din <= x"ffce131d";
		wait for Clk_period;
		Addr <=  "0010010100100";
		Trees_din <= x"002d131d";
		wait for Clk_period;
		Addr <=  "0010010100101";
		Trees_din <= x"00fdce08";
		wait for Clk_period;
		Addr <=  "0010010100110";
		Trees_din <= x"0702a704";
		wait for Clk_period;
		Addr <=  "0010010100111";
		Trees_din <= x"0076131d";
		wait for Clk_period;
		Addr <=  "0010010101000";
		Trees_din <= x"ff7a131d";
		wait for Clk_period;
		Addr <=  "0010010101001";
		Trees_din <= x"12005a04";
		wait for Clk_period;
		Addr <=  "0010010101010";
		Trees_din <= x"ffdf131d";
		wait for Clk_period;
		Addr <=  "0010010101011";
		Trees_din <= x"0098131d";
		wait for Clk_period;
		Addr <=  "0010010101100";
		Trees_din <= x"000e191c";
		wait for Clk_period;
		Addr <=  "0010010101101";
		Trees_din <= x"08002408";
		wait for Clk_period;
		Addr <=  "0010010101110";
		Trees_din <= x"08002204";
		wait for Clk_period;
		Addr <=  "0010010101111";
		Trees_din <= x"005b131d";
		wait for Clk_period;
		Addr <=  "0010010110000";
		Trees_din <= x"ffa3131d";
		wait for Clk_period;
		Addr <=  "0010010110001";
		Trees_din <= x"000bb508";
		wait for Clk_period;
		Addr <=  "0010010110010";
		Trees_din <= x"04f68e04";
		wait for Clk_period;
		Addr <=  "0010010110011";
		Trees_din <= x"0026131d";
		wait for Clk_period;
		Addr <=  "0010010110100";
		Trees_din <= x"009b131d";
		wait for Clk_period;
		Addr <=  "0010010110101";
		Trees_din <= x"03f7a104";
		wait for Clk_period;
		Addr <=  "0010010110110";
		Trees_din <= x"0090131d";
		wait for Clk_period;
		Addr <=  "0010010110111";
		Trees_din <= x"16006f04";
		wait for Clk_period;
		Addr <=  "0010010111000";
		Trees_din <= x"0064131d";
		wait for Clk_period;
		Addr <=  "0010010111001";
		Trees_din <= x"ff2f131d";
		wait for Clk_period;
		Addr <=  "0010010111010";
		Trees_din <= x"0900aa08";
		wait for Clk_period;
		Addr <=  "0010010111011";
		Trees_din <= x"1f028304";
		wait for Clk_period;
		Addr <=  "0010010111100";
		Trees_din <= x"0090131d";
		wait for Clk_period;
		Addr <=  "0010010111101";
		Trees_din <= x"fff5131d";
		wait for Clk_period;
		Addr <=  "0010010111110";
		Trees_din <= x"0113f80c";
		wait for Clk_period;
		Addr <=  "0010010111111";
		Trees_din <= x"0e002504";
		wait for Clk_period;
		Addr <=  "0010011000000";
		Trees_din <= x"0080131d";
		wait for Clk_period;
		Addr <=  "0010011000001";
		Trees_din <= x"02031504";
		wait for Clk_period;
		Addr <=  "0010011000010";
		Trees_din <= x"002b131d";
		wait for Clk_period;
		Addr <=  "0010011000011";
		Trees_din <= x"ff8c131d";
		wait for Clk_period;
		Addr <=  "0010011000100";
		Trees_din <= x"0d013b04";
		wait for Clk_period;
		Addr <=  "0010011000101";
		Trees_din <= x"0087131d";
		wait for Clk_period;
		Addr <=  "0010011000110";
		Trees_din <= x"ffe6131d";
		wait for Clk_period;
		Addr <=  "0010011000111";
		Trees_din <= x"0111b048";
		wait for Clk_period;
		Addr <=  "0010011001000";
		Trees_din <= x"01032f0c";
		wait for Clk_period;
		Addr <=  "0010011001001";
		Trees_din <= x"0c00bb04";
		wait for Clk_period;
		Addr <=  "0010011001010";
		Trees_din <= x"ff741411";
		wait for Clk_period;
		Addr <=  "0010011001011";
		Trees_din <= x"16006004";
		wait for Clk_period;
		Addr <=  "0010011001100";
		Trees_din <= x"ff8e1411";
		wait for Clk_period;
		Addr <=  "0010011001101";
		Trees_din <= x"008c1411";
		wait for Clk_period;
		Addr <=  "0010011001110";
		Trees_din <= x"1402271c";
		wait for Clk_period;
		Addr <=  "0010011001111";
		Trees_din <= x"03f5d50c";
		wait for Clk_period;
		Addr <=  "0010011010000";
		Trees_din <= x"1700bf08";
		wait for Clk_period;
		Addr <=  "0010011010001";
		Trees_din <= x"17f82f04";
		wait for Clk_period;
		Addr <=  "0010011010010";
		Trees_din <= x"004c1411";
		wait for Clk_period;
		Addr <=  "0010011010011";
		Trees_din <= x"ff611411";
		wait for Clk_period;
		Addr <=  "0010011010100";
		Trees_din <= x"00991411";
		wait for Clk_period;
		Addr <=  "0010011010101";
		Trees_din <= x"03fa9508";
		wait for Clk_period;
		Addr <=  "0010011010110";
		Trees_din <= x"0b00b304";
		wait for Clk_period;
		Addr <=  "0010011010111";
		Trees_din <= x"00901411";
		wait for Clk_period;
		Addr <=  "0010011011000";
		Trees_din <= x"ffbd1411";
		wait for Clk_period;
		Addr <=  "0010011011001";
		Trees_din <= x"0006c204";
		wait for Clk_period;
		Addr <=  "0010011011010";
		Trees_din <= x"005b1411";
		wait for Clk_period;
		Addr <=  "0010011011011";
		Trees_din <= x"ff771411";
		wait for Clk_period;
		Addr <=  "0010011011100";
		Trees_din <= x"04020710";
		wait for Clk_period;
		Addr <=  "0010011011101";
		Trees_din <= x"03f47608";
		wait for Clk_period;
		Addr <=  "0010011011110";
		Trees_din <= x"0900e304";
		wait for Clk_period;
		Addr <=  "0010011011111";
		Trees_din <= x"00921411";
		wait for Clk_period;
		Addr <=  "0010011100000";
		Trees_din <= x"ffcc1411";
		wait for Clk_period;
		Addr <=  "0010011100001";
		Trees_din <= x"1f028804";
		wait for Clk_period;
		Addr <=  "0010011100010";
		Trees_din <= x"00001411";
		wait for Clk_period;
		Addr <=  "0010011100011";
		Trees_din <= x"008a1411";
		wait for Clk_period;
		Addr <=  "0010011100100";
		Trees_din <= x"0011e808";
		wait for Clk_period;
		Addr <=  "0010011100101";
		Trees_din <= x"1f028504";
		wait for Clk_period;
		Addr <=  "0010011100110";
		Trees_din <= x"004e1411";
		wait for Clk_period;
		Addr <=  "0010011100111";
		Trees_din <= x"ff6c1411";
		wait for Clk_period;
		Addr <=  "0010011101000";
		Trees_din <= x"10003d04";
		wait for Clk_period;
		Addr <=  "0010011101001";
		Trees_din <= x"003c1411";
		wait for Clk_period;
		Addr <=  "0010011101010";
		Trees_din <= x"ff771411";
		wait for Clk_period;
		Addr <=  "0010011101011";
		Trees_din <= x"000b7d0c";
		wait for Clk_period;
		Addr <=  "0010011101100";
		Trees_din <= x"11000004";
		wait for Clk_period;
		Addr <=  "0010011101101";
		Trees_din <= x"ffe31411";
		wait for Clk_period;
		Addr <=  "0010011101110";
		Trees_din <= x"11032604";
		wait for Clk_period;
		Addr <=  "0010011101111";
		Trees_din <= x"00991411";
		wait for Clk_period;
		Addr <=  "0010011110000";
		Trees_din <= x"00211411";
		wait for Clk_period;
		Addr <=  "0010011110001";
		Trees_din <= x"17f7bc14";
		wait for Clk_period;
		Addr <=  "0010011110010";
		Trees_din <= x"03f7a10c";
		wait for Clk_period;
		Addr <=  "0010011110011";
		Trees_din <= x"01134408";
		wait for Clk_period;
		Addr <=  "0010011110100";
		Trees_din <= x"01125404";
		wait for Clk_period;
		Addr <=  "0010011110101";
		Trees_din <= x"005d1411";
		wait for Clk_period;
		Addr <=  "0010011110110";
		Trees_din <= x"ff961411";
		wait for Clk_period;
		Addr <=  "0010011110111";
		Trees_din <= x"008a1411";
		wait for Clk_period;
		Addr <=  "0010011111000";
		Trees_din <= x"03f82704";
		wait for Clk_period;
		Addr <=  "0010011111001";
		Trees_din <= x"fefb1411";
		wait for Clk_period;
		Addr <=  "0010011111010";
		Trees_din <= x"00211411";
		wait for Clk_period;
		Addr <=  "0010011111011";
		Trees_din <= x"1302e10c";
		wait for Clk_period;
		Addr <=  "0010011111100";
		Trees_din <= x"1302d008";
		wait for Clk_period;
		Addr <=  "0010011111101";
		Trees_din <= x"04012604";
		wait for Clk_period;
		Addr <=  "0010011111110";
		Trees_din <= x"00821411";
		wait for Clk_period;
		Addr <=  "0010011111111";
		Trees_din <= x"ffd91411";
		wait for Clk_period;
		Addr <=  "0010100000000";
		Trees_din <= x"ff481411";
		wait for Clk_period;
		Addr <=  "0010100000001";
		Trees_din <= x"0f000304";
		wait for Clk_period;
		Addr <=  "0010100000010";
		Trees_din <= x"00031411";
		wait for Clk_period;
		Addr <=  "0010100000011";
		Trees_din <= x"00961411";
		wait for Clk_period;
		Addr <=  "0010100000100";
		Trees_din <= x"0111c268";
		wait for Clk_period;
		Addr <=  "0010100000101";
		Trees_din <= x"0109172c";
		wait for Clk_period;
		Addr <=  "0010100000110";
		Trees_din <= x"0a003d0c";
		wait for Clk_period;
		Addr <=  "0010100000111";
		Trees_din <= x"16003f08";
		wait for Clk_period;
		Addr <=  "0010100001000";
		Trees_din <= x"06034b04";
		wait for Clk_period;
		Addr <=  "0010100001001";
		Trees_din <= x"ffea1535";
		wait for Clk_period;
		Addr <=  "0010100001010";
		Trees_din <= x"00801535";
		wait for Clk_period;
		Addr <=  "0010100001011";
		Trees_din <= x"ff601535";
		wait for Clk_period;
		Addr <=  "0010100001100";
		Trees_din <= x"0a004310";
		wait for Clk_period;
		Addr <=  "0010100001101";
		Trees_din <= x"12007708";
		wait for Clk_period;
		Addr <=  "0010100001110";
		Trees_din <= x"15003904";
		wait for Clk_period;
		Addr <=  "0010100001111";
		Trees_din <= x"01051535";
		wait for Clk_period;
		Addr <=  "0010100010000";
		Trees_din <= x"00331535";
		wait for Clk_period;
		Addr <=  "0010100010001";
		Trees_din <= x"0900d904";
		wait for Clk_period;
		Addr <=  "0010100010010";
		Trees_din <= x"00451535";
		wait for Clk_period;
		Addr <=  "0010100010011";
		Trees_din <= x"ff9c1535";
		wait for Clk_period;
		Addr <=  "0010100010100";
		Trees_din <= x"03f8e608";
		wait for Clk_period;
		Addr <=  "0010100010101";
		Trees_din <= x"0f000704";
		wait for Clk_period;
		Addr <=  "0010100010110";
		Trees_din <= x"00401535";
		wait for Clk_period;
		Addr <=  "0010100010111";
		Trees_din <= x"ffb11535";
		wait for Clk_period;
		Addr <=  "0010100011000";
		Trees_din <= x"05f77a04";
		wait for Clk_period;
		Addr <=  "0010100011001";
		Trees_din <= x"ff5b1535";
		wait for Clk_period;
		Addr <=  "0010100011010";
		Trees_din <= x"ffe81535";
		wait for Clk_period;
		Addr <=  "0010100011011";
		Trees_din <= x"1402ee1c";
		wait for Clk_period;
		Addr <=  "0010100011100";
		Trees_din <= x"10004e10";
		wait for Clk_period;
		Addr <=  "0010100011101";
		Trees_din <= x"19000108";
		wait for Clk_period;
		Addr <=  "0010100011110";
		Trees_din <= x"08004704";
		wait for Clk_period;
		Addr <=  "0010100011111";
		Trees_din <= x"00c81535";
		wait for Clk_period;
		Addr <=  "0010100100000";
		Trees_din <= x"fff11535";
		wait for Clk_period;
		Addr <=  "0010100100001";
		Trees_din <= x"19000204";
		wait for Clk_period;
		Addr <=  "0010100100010";
		Trees_din <= x"ff4b1535";
		wait for Clk_period;
		Addr <=  "0010100100011";
		Trees_din <= x"00401535";
		wait for Clk_period;
		Addr <=  "0010100100100";
		Trees_din <= x"0600a108";
		wait for Clk_period;
		Addr <=  "0010100100101";
		Trees_din <= x"1b027e04";
		wait for Clk_period;
		Addr <=  "0010100100110";
		Trees_din <= x"ff401535";
		wait for Clk_period;
		Addr <=  "0010100100111";
		Trees_din <= x"00041535";
		wait for Clk_period;
		Addr <=  "0010100101000";
		Trees_din <= x"00841535";
		wait for Clk_period;
		Addr <=  "0010100101001";
		Trees_din <= x"1afadd10";
		wait for Clk_period;
		Addr <=  "0010100101010";
		Trees_din <= x"1e028308";
		wait for Clk_period;
		Addr <=  "0010100101011";
		Trees_din <= x"0a003e04";
		wait for Clk_period;
		Addr <=  "0010100101100";
		Trees_din <= x"00261535";
		wait for Clk_period;
		Addr <=  "0010100101101";
		Trees_din <= x"ff4a1535";
		wait for Clk_period;
		Addr <=  "0010100101110";
		Trees_din <= x"0d001c04";
		wait for Clk_period;
		Addr <=  "0010100101111";
		Trees_din <= x"ffad1535";
		wait for Clk_period;
		Addr <=  "0010100110000";
		Trees_din <= x"00391535";
		wait for Clk_period;
		Addr <=  "0010100110001";
		Trees_din <= x"15003608";
		wait for Clk_period;
		Addr <=  "0010100110010";
		Trees_din <= x"06ff0e04";
		wait for Clk_period;
		Addr <=  "0010100110011";
		Trees_din <= x"ffff1535";
		wait for Clk_period;
		Addr <=  "0010100110100";
		Trees_din <= x"007a1535";
		wait for Clk_period;
		Addr <=  "0010100110101";
		Trees_din <= x"16006204";
		wait for Clk_period;
		Addr <=  "0010100110110";
		Trees_din <= x"ffc01535";
		wait for Clk_period;
		Addr <=  "0010100110111";
		Trees_din <= x"00121535";
		wait for Clk_period;
		Addr <=  "0010100111000";
		Trees_din <= x"000b7d0c";
		wait for Clk_period;
		Addr <=  "0010100111001";
		Trees_din <= x"11000004";
		wait for Clk_period;
		Addr <=  "0010100111010";
		Trees_din <= x"ffe11535";
		wait for Clk_period;
		Addr <=  "0010100111011";
		Trees_din <= x"11032604";
		wait for Clk_period;
		Addr <=  "0010100111100";
		Trees_din <= x"00971535";
		wait for Clk_period;
		Addr <=  "0010100111101";
		Trees_din <= x"001e1535";
		wait for Clk_period;
		Addr <=  "0010100111110";
		Trees_din <= x"03f7a110";
		wait for Clk_period;
		Addr <=  "0010100111111";
		Trees_din <= x"0a00480c";
		wait for Clk_period;
		Addr <=  "0010101000000";
		Trees_din <= x"0a004708";
		wait for Clk_period;
		Addr <=  "0010101000001";
		Trees_din <= x"19000004";
		wait for Clk_period;
		Addr <=  "0010101000010";
		Trees_din <= x"00131535";
		wait for Clk_period;
		Addr <=  "0010101000011";
		Trees_din <= x"008f1535";
		wait for Clk_period;
		Addr <=  "0010101000100";
		Trees_din <= x"ff781535";
		wait for Clk_period;
		Addr <=  "0010101000101";
		Trees_din <= x"008a1535";
		wait for Clk_period;
		Addr <=  "0010101000110";
		Trees_din <= x"03f82708";
		wait for Clk_period;
		Addr <=  "0010101000111";
		Trees_din <= x"0900d504";
		wait for Clk_period;
		Addr <=  "0010101001000";
		Trees_din <= x"ffb71535";
		wait for Clk_period;
		Addr <=  "0010101001001";
		Trees_din <= x"ff011535";
		wait for Clk_period;
		Addr <=  "0010101001010";
		Trees_din <= x"1c026204";
		wait for Clk_period;
		Addr <=  "0010101001011";
		Trees_din <= x"00191535";
		wait for Clk_period;
		Addr <=  "0010101001100";
		Trees_din <= x"00731535";
		wait for Clk_period;
		Addr <=  "0010101001101";
		Trees_din <= x"0111c23c";
		wait for Clk_period;
		Addr <=  "0010101001110";
		Trees_din <= x"01032f0c";
		wait for Clk_period;
		Addr <=  "0010101001111";
		Trees_din <= x"0c00bb04";
		wait for Clk_period;
		Addr <=  "0010101010000";
		Trees_din <= x"ff771611";
		wait for Clk_period;
		Addr <=  "0010101010001";
		Trees_din <= x"16006004";
		wait for Clk_period;
		Addr <=  "0010101010010";
		Trees_din <= x"ff941611";
		wait for Clk_period;
		Addr <=  "0010101010011";
		Trees_din <= x"00731611";
		wait for Clk_period;
		Addr <=  "0010101010100";
		Trees_din <= x"1600a720";
		wait for Clk_period;
		Addr <=  "0010101010101";
		Trees_din <= x"10005610";
		wait for Clk_period;
		Addr <=  "0010101010110";
		Trees_din <= x"16009608";
		wait for Clk_period;
		Addr <=  "0010101010111";
		Trees_din <= x"15004c04";
		wait for Clk_period;
		Addr <=  "0010101011000";
		Trees_din <= x"000d1611";
		wait for Clk_period;
		Addr <=  "0010101011001";
		Trees_din <= x"ffad1611";
		wait for Clk_period;
		Addr <=  "0010101011010";
		Trees_din <= x"02019d04";
		wait for Clk_period;
		Addr <=  "0010101011011";
		Trees_din <= x"ffd11611";
		wait for Clk_period;
		Addr <=  "0010101011100";
		Trees_din <= x"00ba1611";
		wait for Clk_period;
		Addr <=  "0010101011101";
		Trees_din <= x"1b026c08";
		wait for Clk_period;
		Addr <=  "0010101011110";
		Trees_din <= x"05f4f804";
		wait for Clk_period;
		Addr <=  "0010101011111";
		Trees_din <= x"ffe91611";
		wait for Clk_period;
		Addr <=  "0010101100000";
		Trees_din <= x"ff521611";
		wait for Clk_period;
		Addr <=  "0010101100001";
		Trees_din <= x"010ae204";
		wait for Clk_period;
		Addr <=  "0010101100010";
		Trees_din <= x"ff871611";
		wait for Clk_period;
		Addr <=  "0010101100011";
		Trees_din <= x"006b1611";
		wait for Clk_period;
		Addr <=  "0010101100100";
		Trees_din <= x"0900d908";
		wait for Clk_period;
		Addr <=  "0010101100101";
		Trees_din <= x"08004504";
		wait for Clk_period;
		Addr <=  "0010101100110";
		Trees_din <= x"00a61611";
		wait for Clk_period;
		Addr <=  "0010101100111";
		Trees_din <= x"ffff1611";
		wait for Clk_period;
		Addr <=  "0010101101000";
		Trees_din <= x"010d9f04";
		wait for Clk_period;
		Addr <=  "0010101101001";
		Trees_din <= x"ff751611";
		wait for Clk_period;
		Addr <=  "0010101101010";
		Trees_din <= x"004e1611";
		wait for Clk_period;
		Addr <=  "0010101101011";
		Trees_din <= x"000b7d0c";
		wait for Clk_period;
		Addr <=  "0010101101100";
		Trees_din <= x"11000004";
		wait for Clk_period;
		Addr <=  "0010101101101";
		Trees_din <= x"ffe41611";
		wait for Clk_period;
		Addr <=  "0010101101110";
		Trees_din <= x"16009104";
		wait for Clk_period;
		Addr <=  "0010101101111";
		Trees_din <= x"00941611";
		wait for Clk_period;
		Addr <=  "0010101110000";
		Trees_din <= x"00201611";
		wait for Clk_period;
		Addr <=  "0010101110001";
		Trees_din <= x"17f7bc14";
		wait for Clk_period;
		Addr <=  "0010101110010";
		Trees_din <= x"03f7a10c";
		wait for Clk_period;
		Addr <=  "0010101110011";
		Trees_din <= x"01134408";
		wait for Clk_period;
		Addr <=  "0010101110100";
		Trees_din <= x"01125404";
		wait for Clk_period;
		Addr <=  "0010101110101";
		Trees_din <= x"00741611";
		wait for Clk_period;
		Addr <=  "0010101110110";
		Trees_din <= x"ff981611";
		wait for Clk_period;
		Addr <=  "0010101110111";
		Trees_din <= x"00801611";
		wait for Clk_period;
		Addr <=  "0010101111000";
		Trees_din <= x"03f82704";
		wait for Clk_period;
		Addr <=  "0010101111001";
		Trees_din <= x"ff261611";
		wait for Clk_period;
		Addr <=  "0010101111010";
		Trees_din <= x"00141611";
		wait for Clk_period;
		Addr <=  "0010101111011";
		Trees_din <= x"0f009408";
		wait for Clk_period;
		Addr <=  "0010101111100";
		Trees_din <= x"1403ff04";
		wait for Clk_period;
		Addr <=  "0010101111101";
		Trees_din <= x"008d1611";
		wait for Clk_period;
		Addr <=  "0010101111110";
		Trees_din <= x"00081611";
		wait for Clk_period;
		Addr <=  "0010101111111";
		Trees_din <= x"1302e108";
		wait for Clk_period;
		Addr <=  "0010110000000";
		Trees_din <= x"1302cb04";
		wait for Clk_period;
		Addr <=  "0010110000001";
		Trees_din <= x"00261611";
		wait for Clk_period;
		Addr <=  "0010110000010";
		Trees_din <= x"ff5d1611";
		wait for Clk_period;
		Addr <=  "0010110000011";
		Trees_din <= x"00701611";
		wait for Clk_period;
		Addr <=  "0010110000100";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0010110000101";
		Trees_din <= x"0111c264";
		wait for Clk_period;
		Addr <=  "0010110000110";
		Trees_din <= x"01054b24";
		wait for Clk_period;
		Addr <=  "0010110000111";
		Trees_din <= x"15003914";
		wait for Clk_period;
		Addr <=  "0010110001000";
		Trees_din <= x"11017c10";
		wait for Clk_period;
		Addr <=  "0010110001001";
		Trees_din <= x"00054f08";
		wait for Clk_period;
		Addr <=  "0010110001010";
		Trees_din <= x"0002aa04";
		wait for Clk_period;
		Addr <=  "0010110001011";
		Trees_din <= x"00141739";
		wait for Clk_period;
		Addr <=  "0010110001100";
		Trees_din <= x"00d91739";
		wait for Clk_period;
		Addr <=  "0010110001101";
		Trees_din <= x"1f026204";
		wait for Clk_period;
		Addr <=  "0010110001110";
		Trees_din <= x"00121739";
		wait for Clk_period;
		Addr <=  "0010110001111";
		Trees_din <= x"ff971739";
		wait for Clk_period;
		Addr <=  "0010110010000";
		Trees_din <= x"ff881739";
		wait for Clk_period;
		Addr <=  "0010110010001";
		Trees_din <= x"0900e404";
		wait for Clk_period;
		Addr <=  "0010110010010";
		Trees_din <= x"ff6e1739";
		wait for Clk_period;
		Addr <=  "0010110010011";
		Trees_din <= x"0900e504";
		wait for Clk_period;
		Addr <=  "0010110010100";
		Trees_din <= x"00881739";
		wait for Clk_period;
		Addr <=  "0010110010101";
		Trees_din <= x"0002aa04";
		wait for Clk_period;
		Addr <=  "0010110010110";
		Trees_din <= x"000a1739";
		wait for Clk_period;
		Addr <=  "0010110010111";
		Trees_din <= x"ff831739";
		wait for Clk_period;
		Addr <=  "0010110011000";
		Trees_din <= x"04020720";
		wait for Clk_period;
		Addr <=  "0010110011001";
		Trees_din <= x"03f47610";
		wait for Clk_period;
		Addr <=  "0010110011010";
		Trees_din <= x"0b008608";
		wait for Clk_period;
		Addr <=  "0010110011011";
		Trees_din <= x"07f9f604";
		wait for Clk_period;
		Addr <=  "0010110011100";
		Trees_din <= x"001f1739";
		wait for Clk_period;
		Addr <=  "0010110011101";
		Trees_din <= x"00b31739";
		wait for Clk_period;
		Addr <=  "0010110011110";
		Trees_din <= x"12009004";
		wait for Clk_period;
		Addr <=  "0010110011111";
		Trees_din <= x"ff601739";
		wait for Clk_period;
		Addr <=  "0010110100000";
		Trees_din <= x"00371739";
		wait for Clk_period;
		Addr <=  "0010110100001";
		Trees_din <= x"03f4de08";
		wait for Clk_period;
		Addr <=  "0010110100010";
		Trees_din <= x"04010f04";
		wait for Clk_period;
		Addr <=  "0010110100011";
		Trees_din <= x"ff5e1739";
		wait for Clk_period;
		Addr <=  "0010110100100";
		Trees_din <= x"00761739";
		wait for Clk_period;
		Addr <=  "0010110100101";
		Trees_din <= x"0401d104";
		wait for Clk_period;
		Addr <=  "0010110100110";
		Trees_din <= x"00061739";
		wait for Clk_period;
		Addr <=  "0010110100111";
		Trees_din <= x"ff791739";
		wait for Clk_period;
		Addr <=  "0010110101000";
		Trees_din <= x"0900e610";
		wait for Clk_period;
		Addr <=  "0010110101001";
		Trees_din <= x"010b1308";
		wait for Clk_period;
		Addr <=  "0010110101010";
		Trees_din <= x"16004d04";
		wait for Clk_period;
		Addr <=  "0010110101011";
		Trees_din <= x"008e1739";
		wait for Clk_period;
		Addr <=  "0010110101100";
		Trees_din <= x"ffa01739";
		wait for Clk_period;
		Addr <=  "0010110101101";
		Trees_din <= x"12008404";
		wait for Clk_period;
		Addr <=  "0010110101110";
		Trees_din <= x"005c1739";
		wait for Clk_period;
		Addr <=  "0010110101111";
		Trees_din <= x"ffbe1739";
		wait for Clk_period;
		Addr <=  "0010110110000";
		Trees_din <= x"0c009408";
		wait for Clk_period;
		Addr <=  "0010110110001";
		Trees_din <= x"07f59c04";
		wait for Clk_period;
		Addr <=  "0010110110010";
		Trees_din <= x"00441739";
		wait for Clk_period;
		Addr <=  "0010110110011";
		Trees_din <= x"ff8c1739";
		wait for Clk_period;
		Addr <=  "0010110110100";
		Trees_din <= x"12006f04";
		wait for Clk_period;
		Addr <=  "0010110110101";
		Trees_din <= x"01241739";
		wait for Clk_period;
		Addr <=  "0010110110110";
		Trees_din <= x"00681739";
		wait for Clk_period;
		Addr <=  "0010110110111";
		Trees_din <= x"000b7d0c";
		wait for Clk_period;
		Addr <=  "0010110111000";
		Trees_din <= x"21001408";
		wait for Clk_period;
		Addr <=  "0010110111001";
		Trees_din <= x"16009104";
		wait for Clk_period;
		Addr <=  "0010110111010";
		Trees_din <= x"00921739";
		wait for Clk_period;
		Addr <=  "0010110111011";
		Trees_din <= x"001f1739";
		wait for Clk_period;
		Addr <=  "0010110111100";
		Trees_din <= x"ffdc1739";
		wait for Clk_period;
		Addr <=  "0010110111101";
		Trees_din <= x"08003f14";
		wait for Clk_period;
		Addr <=  "0010110111110";
		Trees_din <= x"0d00a60c";
		wait for Clk_period;
		Addr <=  "0010110111111";
		Trees_din <= x"18002508";
		wait for Clk_period;
		Addr <=  "0010111000000";
		Trees_din <= x"01130b04";
		wait for Clk_period;
		Addr <=  "0010111000001";
		Trees_din <= x"ffab1739";
		wait for Clk_period;
		Addr <=  "0010111000010";
		Trees_din <= x"00671739";
		wait for Clk_period;
		Addr <=  "0010111000011";
		Trees_din <= x"007d1739";
		wait for Clk_period;
		Addr <=  "0010111000100";
		Trees_din <= x"1101af04";
		wait for Clk_period;
		Addr <=  "0010111000101";
		Trees_din <= x"ff3b1739";
		wait for Clk_period;
		Addr <=  "0010111000110";
		Trees_din <= x"001b1739";
		wait for Clk_period;
		Addr <=  "0010111000111";
		Trees_din <= x"03f5180c";
		wait for Clk_period;
		Addr <=  "0010111001000";
		Trees_din <= x"0b007008";
		wait for Clk_period;
		Addr <=  "0010111001001";
		Trees_din <= x"0b006c04";
		wait for Clk_period;
		Addr <=  "0010111001010";
		Trees_din <= x"001a1739";
		wait for Clk_period;
		Addr <=  "0010111001011";
		Trees_din <= x"ff8e1739";
		wait for Clk_period;
		Addr <=  "0010111001100";
		Trees_din <= x"00691739";
		wait for Clk_period;
		Addr <=  "0010111001101";
		Trees_din <= x"00841739";
		wait for Clk_period;
		Addr <=  "0010111001110";
		Trees_din <= x"0111f870";
		wait for Clk_period;
		Addr <=  "0010111001111";
		Trees_din <= x"06ff2534";
		wait for Clk_period;
		Addr <=  "0010111010000";
		Trees_din <= x"10005c20";
		wait for Clk_period;
		Addr <=  "0010111010001";
		Trees_din <= x"010fcb10";
		wait for Clk_period;
		Addr <=  "0010111010010";
		Trees_din <= x"15004a08";
		wait for Clk_period;
		Addr <=  "0010111010011";
		Trees_din <= x"0e002804";
		wait for Clk_period;
		Addr <=  "0010111010100";
		Trees_din <= x"ffd11875";
		wait for Clk_period;
		Addr <=  "0010111010101";
		Trees_din <= x"00061875";
		wait for Clk_period;
		Addr <=  "0010111010110";
		Trees_din <= x"0900ea04";
		wait for Clk_period;
		Addr <=  "0010111010111";
		Trees_din <= x"ff7a1875";
		wait for Clk_period;
		Addr <=  "0010111011000";
		Trees_din <= x"00ac1875";
		wait for Clk_period;
		Addr <=  "0010111011001";
		Trees_din <= x"0f000008";
		wait for Clk_period;
		Addr <=  "0010111011010";
		Trees_din <= x"11000904";
		wait for Clk_period;
		Addr <=  "0010111011011";
		Trees_din <= x"004d1875";
		wait for Clk_period;
		Addr <=  "0010111011100";
		Trees_din <= x"ff5f1875";
		wait for Clk_period;
		Addr <=  "0010111011101";
		Trees_din <= x"0f000404";
		wait for Clk_period;
		Addr <=  "0010111011110";
		Trees_din <= x"009b1875";
		wait for Clk_period;
		Addr <=  "0010111011111";
		Trees_din <= x"001c1875";
		wait for Clk_period;
		Addr <=  "0010111100000";
		Trees_din <= x"0a00520c";
		wait for Clk_period;
		Addr <=  "0010111100001";
		Trees_din <= x"06fc9a04";
		wait for Clk_period;
		Addr <=  "0010111100010";
		Trees_din <= x"006e1875";
		wait for Clk_period;
		Addr <=  "0010111100011";
		Trees_din <= x"0f000004";
		wait for Clk_period;
		Addr <=  "0010111100100";
		Trees_din <= x"ff8e1875";
		wait for Clk_period;
		Addr <=  "0010111100101";
		Trees_din <= x"001b1875";
		wait for Clk_period;
		Addr <=  "0010111100110";
		Trees_din <= x"08003c04";
		wait for Clk_period;
		Addr <=  "0010111100111";
		Trees_din <= x"00b81875";
		wait for Clk_period;
		Addr <=  "0010111101000";
		Trees_din <= x"001f1875";
		wait for Clk_period;
		Addr <=  "0010111101001";
		Trees_din <= x"0a003d20";
		wait for Clk_period;
		Addr <=  "0010111101010";
		Trees_din <= x"010d0210";
		wait for Clk_period;
		Addr <=  "0010111101011";
		Trees_din <= x"17f9ad08";
		wait for Clk_period;
		Addr <=  "0010111101100";
		Trees_din <= x"02026504";
		wait for Clk_period;
		Addr <=  "0010111101101";
		Trees_din <= x"00451875";
		wait for Clk_period;
		Addr <=  "0010111101110";
		Trees_din <= x"ff631875";
		wait for Clk_period;
		Addr <=  "0010111101111";
		Trees_din <= x"1101a104";
		wait for Clk_period;
		Addr <=  "0010111110000";
		Trees_din <= x"00891875";
		wait for Clk_period;
		Addr <=  "0010111110001";
		Trees_din <= x"ff8d1875";
		wait for Clk_period;
		Addr <=  "0010111110010";
		Trees_din <= x"0b006208";
		wait for Clk_period;
		Addr <=  "0010111110011";
		Trees_din <= x"02048e04";
		wait for Clk_period;
		Addr <=  "0010111110100";
		Trees_din <= x"ff0f1875";
		wait for Clk_period;
		Addr <=  "0010111110101";
		Trees_din <= x"001b1875";
		wait for Clk_period;
		Addr <=  "0010111110110";
		Trees_din <= x"07f93f04";
		wait for Clk_period;
		Addr <=  "0010111110111";
		Trees_din <= x"001f1875";
		wait for Clk_period;
		Addr <=  "0010111111000";
		Trees_din <= x"009e1875";
		wait for Clk_period;
		Addr <=  "0010111111001";
		Trees_din <= x"0b005f0c";
		wait for Clk_period;
		Addr <=  "0010111111010";
		Trees_din <= x"15004504";
		wait for Clk_period;
		Addr <=  "0010111111011";
		Trees_din <= x"ff8d1875";
		wait for Clk_period;
		Addr <=  "0010111111100";
		Trees_din <= x"08004604";
		wait for Clk_period;
		Addr <=  "0010111111101";
		Trees_din <= x"00941875";
		wait for Clk_period;
		Addr <=  "0010111111110";
		Trees_din <= x"ff991875";
		wait for Clk_period;
		Addr <=  "0010111111111";
		Trees_din <= x"16008108";
		wait for Clk_period;
		Addr <=  "0011000000000";
		Trees_din <= x"04ffb204";
		wait for Clk_period;
		Addr <=  "0011000000001";
		Trees_din <= x"00341875";
		wait for Clk_period;
		Addr <=  "0011000000010";
		Trees_din <= x"ffff1875";
		wait for Clk_period;
		Addr <=  "0011000000011";
		Trees_din <= x"0900bf04";
		wait for Clk_period;
		Addr <=  "0011000000100";
		Trees_din <= x"fff11875";
		wait for Clk_period;
		Addr <=  "0011000000101";
		Trees_din <= x"ff731875";
		wait for Clk_period;
		Addr <=  "0011000000110";
		Trees_din <= x"000e1910";
		wait for Clk_period;
		Addr <=  "0011000000111";
		Trees_din <= x"08003008";
		wait for Clk_period;
		Addr <=  "0011000001000";
		Trees_din <= x"0900c804";
		wait for Clk_period;
		Addr <=  "0011000001001";
		Trees_din <= x"ffa61875";
		wait for Clk_period;
		Addr <=  "0011000001010";
		Trees_din <= x"00611875";
		wait for Clk_period;
		Addr <=  "0011000001011";
		Trees_din <= x"00013504";
		wait for Clk_period;
		Addr <=  "0011000001100";
		Trees_din <= x"00211875";
		wait for Clk_period;
		Addr <=  "0011000001101";
		Trees_din <= x"00911875";
		wait for Clk_period;
		Addr <=  "0011000001110";
		Trees_din <= x"19000014";
		wait for Clk_period;
		Addr <=  "0011000001111";
		Trees_din <= x"0113880c";
		wait for Clk_period;
		Addr <=  "0011000010000";
		Trees_din <= x"0a004808";
		wait for Clk_period;
		Addr <=  "0011000010001";
		Trees_din <= x"07f81804";
		wait for Clk_period;
		Addr <=  "0011000010010";
		Trees_din <= x"ff711875";
		wait for Clk_period;
		Addr <=  "0011000010011";
		Trees_din <= x"fff21875";
		wait for Clk_period;
		Addr <=  "0011000010100";
		Trees_din <= x"00331875";
		wait for Clk_period;
		Addr <=  "0011000010101";
		Trees_din <= x"0c00b004";
		wait for Clk_period;
		Addr <=  "0011000010110";
		Trees_din <= x"00681875";
		wait for Clk_period;
		Addr <=  "0011000010111";
		Trees_din <= x"00001875";
		wait for Clk_period;
		Addr <=  "0011000011000";
		Trees_din <= x"000f3608";
		wait for Clk_period;
		Addr <=  "0011000011001";
		Trees_din <= x"1f027304";
		wait for Clk_period;
		Addr <=  "0011000011010";
		Trees_din <= x"fffc1875";
		wait for Clk_period;
		Addr <=  "0011000011011";
		Trees_din <= x"000c1875";
		wait for Clk_period;
		Addr <=  "0011000011100";
		Trees_din <= x"00791875";
		wait for Clk_period;
		Addr <=  "0011000011101";
		Trees_din <= x"05f51e64";
		wait for Clk_period;
		Addr <=  "0011000011110";
		Trees_din <= x"03f99440";
		wait for Clk_period;
		Addr <=  "0011000011111";
		Trees_din <= x"04006320";
		wait for Clk_period;
		Addr <=  "0011000100000";
		Trees_din <= x"12007f10";
		wait for Clk_period;
		Addr <=  "0011000100001";
		Trees_din <= x"1b023d08";
		wait for Clk_period;
		Addr <=  "0011000100010";
		Trees_din <= x"05f21d04";
		wait for Clk_period;
		Addr <=  "0011000100011";
		Trees_din <= x"ffef1a01";
		wait for Clk_period;
		Addr <=  "0011000100100";
		Trees_din <= x"00a01a01";
		wait for Clk_period;
		Addr <=  "0011000100101";
		Trees_din <= x"0900e204";
		wait for Clk_period;
		Addr <=  "0011000100110";
		Trees_din <= x"ffc01a01";
		wait for Clk_period;
		Addr <=  "0011000100111";
		Trees_din <= x"00071a01";
		wait for Clk_period;
		Addr <=  "0011000101000";
		Trees_din <= x"0a003f08";
		wait for Clk_period;
		Addr <=  "0011000101001";
		Trees_din <= x"12008b04";
		wait for Clk_period;
		Addr <=  "0011000101010";
		Trees_din <= x"ff671a01";
		wait for Clk_period;
		Addr <=  "0011000101011";
		Trees_din <= x"00531a01";
		wait for Clk_period;
		Addr <=  "0011000101100";
		Trees_din <= x"0b007904";
		wait for Clk_period;
		Addr <=  "0011000101101";
		Trees_din <= x"00cf1a01";
		wait for Clk_period;
		Addr <=  "0011000101110";
		Trees_din <= x"00271a01";
		wait for Clk_period;
		Addr <=  "0011000101111";
		Trees_din <= x"0d002710";
		wait for Clk_period;
		Addr <=  "0011000110000";
		Trees_din <= x"000f5408";
		wait for Clk_period;
		Addr <=  "0011000110001";
		Trees_din <= x"03f8d704";
		wait for Clk_period;
		Addr <=  "0011000110010";
		Trees_din <= x"00a21a01";
		wait for Clk_period;
		Addr <=  "0011000110011";
		Trees_din <= x"ffb61a01";
		wait for Clk_period;
		Addr <=  "0011000110100";
		Trees_din <= x"0f000b04";
		wait for Clk_period;
		Addr <=  "0011000110101";
		Trees_din <= x"ffa41a01";
		wait for Clk_period;
		Addr <=  "0011000110110";
		Trees_din <= x"00761a01";
		wait for Clk_period;
		Addr <=  "0011000110111";
		Trees_din <= x"0900e008";
		wait for Clk_period;
		Addr <=  "0011000111000";
		Trees_din <= x"0a004304";
		wait for Clk_period;
		Addr <=  "0011000111001";
		Trees_din <= x"00731a01";
		wait for Clk_period;
		Addr <=  "0011000111010";
		Trees_din <= x"ffee1a01";
		wait for Clk_period;
		Addr <=  "0011000111011";
		Trees_din <= x"07f89204";
		wait for Clk_period;
		Addr <=  "0011000111100";
		Trees_din <= x"00151a01";
		wait for Clk_period;
		Addr <=  "0011000111101";
		Trees_din <= x"ff721a01";
		wait for Clk_period;
		Addr <=  "0011000111110";
		Trees_din <= x"04fed714";
		wait for Clk_period;
		Addr <=  "0011000111111";
		Trees_din <= x"0208ef10";
		wait for Clk_period;
		Addr <=  "0011001000000";
		Trees_din <= x"0900d908";
		wait for Clk_period;
		Addr <=  "0011001000001";
		Trees_din <= x"04fc2904";
		wait for Clk_period;
		Addr <=  "0011001000010";
		Trees_din <= x"004f1a01";
		wait for Clk_period;
		Addr <=  "0011001000011";
		Trees_din <= x"ffbb1a01";
		wait for Clk_period;
		Addr <=  "0011001000100";
		Trees_din <= x"0203e904";
		wait for Clk_period;
		Addr <=  "0011001000101";
		Trees_din <= x"fff11a01";
		wait for Clk_period;
		Addr <=  "0011001000110";
		Trees_din <= x"009a1a01";
		wait for Clk_period;
		Addr <=  "0011001000111";
		Trees_din <= x"ff6c1a01";
		wait for Clk_period;
		Addr <=  "0011001001000";
		Trees_din <= x"17f72504";
		wait for Clk_period;
		Addr <=  "0011001001001";
		Trees_din <= x"ffbb1a01";
		wait for Clk_period;
		Addr <=  "0011001001010";
		Trees_din <= x"0602d008";
		wait for Clk_period;
		Addr <=  "0011001001011";
		Trees_din <= x"0a004704";
		wait for Clk_period;
		Addr <=  "0011001001100";
		Trees_din <= x"00f71a01";
		wait for Clk_period;
		Addr <=  "0011001001101";
		Trees_din <= x"005f1a01";
		wait for Clk_period;
		Addr <=  "0011001001110";
		Trees_din <= x"ffbe1a01";
		wait for Clk_period;
		Addr <=  "0011001001111";
		Trees_din <= x"02044d38";
		wait for Clk_period;
		Addr <=  "0011001010000";
		Trees_din <= x"010ab118";
		wait for Clk_period;
		Addr <=  "0011001010001";
		Trees_din <= x"1d02840c";
		wait for Clk_period;
		Addr <=  "0011001010010";
		Trees_din <= x"0008fe08";
		wait for Clk_period;
		Addr <=  "0011001010011";
		Trees_din <= x"06fd5904";
		wait for Clk_period;
		Addr <=  "0011001010100";
		Trees_din <= x"ff901a01";
		wait for Clk_period;
		Addr <=  "0011001010101";
		Trees_din <= x"00111a01";
		wait for Clk_period;
		Addr <=  "0011001010110";
		Trees_din <= x"ff691a01";
		wait for Clk_period;
		Addr <=  "0011001010111";
		Trees_din <= x"12007804";
		wait for Clk_period;
		Addr <=  "0011001011000";
		Trees_din <= x"ffde1a01";
		wait for Clk_period;
		Addr <=  "0011001011001";
		Trees_din <= x"03f7f604";
		wait for Clk_period;
		Addr <=  "0011001011010";
		Trees_din <= x"00eb1a01";
		wait for Clk_period;
		Addr <=  "0011001011011";
		Trees_din <= x"00091a01";
		wait for Clk_period;
		Addr <=  "0011001011100";
		Trees_din <= x"06febc10";
		wait for Clk_period;
		Addr <=  "0011001011101";
		Trees_din <= x"1801ca08";
		wait for Clk_period;
		Addr <=  "0011001011110";
		Trees_din <= x"18018d04";
		wait for Clk_period;
		Addr <=  "0011001011111";
		Trees_din <= x"000b1a01";
		wait for Clk_period;
		Addr <=  "0011001100000";
		Trees_din <= x"ff081a01";
		wait for Clk_period;
		Addr <=  "0011001100001";
		Trees_din <= x"11029e04";
		wait for Clk_period;
		Addr <=  "0011001100010";
		Trees_din <= x"00b51a01";
		wait for Clk_period;
		Addr <=  "0011001100011";
		Trees_din <= x"00301a01";
		wait for Clk_period;
		Addr <=  "0011001100100";
		Trees_din <= x"18006908";
		wait for Clk_period;
		Addr <=  "0011001100101";
		Trees_din <= x"12006304";
		wait for Clk_period;
		Addr <=  "0011001100110";
		Trees_din <= x"002d1a01";
		wait for Clk_period;
		Addr <=  "0011001100111";
		Trees_din <= x"00bf1a01";
		wait for Clk_period;
		Addr <=  "0011001101000";
		Trees_din <= x"010ae204";
		wait for Clk_period;
		Addr <=  "0011001101001";
		Trees_din <= x"ff5f1a01";
		wait for Clk_period;
		Addr <=  "0011001101010";
		Trees_din <= x"005c1a01";
		wait for Clk_period;
		Addr <=  "0011001101011";
		Trees_din <= x"0a003c0c";
		wait for Clk_period;
		Addr <=  "0011001101100";
		Trees_din <= x"010d5f08";
		wait for Clk_period;
		Addr <=  "0011001101101";
		Trees_din <= x"0a003704";
		wait for Clk_period;
		Addr <=  "0011001101110";
		Trees_din <= x"00011a01";
		wait for Clk_period;
		Addr <=  "0011001101111";
		Trees_din <= x"ff331a01";
		wait for Clk_period;
		Addr <=  "0011001110000";
		Trees_din <= x"00651a01";
		wait for Clk_period;
		Addr <=  "0011001110001";
		Trees_din <= x"0009cb10";
		wait for Clk_period;
		Addr <=  "0011001110010";
		Trees_din <= x"020ce808";
		wait for Clk_period;
		Addr <=  "0011001110011";
		Trees_din <= x"0006b204";
		wait for Clk_period;
		Addr <=  "0011001110100";
		Trees_din <= x"ffe21a01";
		wait for Clk_period;
		Addr <=  "0011001110101";
		Trees_din <= x"00201a01";
		wait for Clk_period;
		Addr <=  "0011001110110";
		Trees_din <= x"07fb5f04";
		wait for Clk_period;
		Addr <=  "0011001110111";
		Trees_din <= x"fff51a01";
		wait for Clk_period;
		Addr <=  "0011001111000";
		Trees_din <= x"01411a01";
		wait for Clk_period;
		Addr <=  "0011001111001";
		Trees_din <= x"0f000008";
		wait for Clk_period;
		Addr <=  "0011001111010";
		Trees_din <= x"06011904";
		wait for Clk_period;
		Addr <=  "0011001111011";
		Trees_din <= x"ff201a01";
		wait for Clk_period;
		Addr <=  "0011001111100";
		Trees_din <= x"00291a01";
		wait for Clk_period;
		Addr <=  "0011001111101";
		Trees_din <= x"08003804";
		wait for Clk_period;
		Addr <=  "0011001111110";
		Trees_din <= x"ff7b1a01";
		wait for Clk_period;
		Addr <=  "0011001111111";
		Trees_din <= x"fffe1a01";
		wait for Clk_period;
		Addr <=  "0011010000000";
		Trees_din <= x"0d009168";
		wait for Clk_period;
		Addr <=  "0011010000001";
		Trees_din <= x"05f3fd38";
		wait for Clk_period;
		Addr <=  "0011010000010";
		Trees_din <= x"11008c20";
		wait for Clk_period;
		Addr <=  "0011010000011";
		Trees_din <= x"1b026e10";
		wait for Clk_period;
		Addr <=  "0011010000100";
		Trees_din <= x"0f001108";
		wait for Clk_period;
		Addr <=  "0011010000101";
		Trees_din <= x"0f000604";
		wait for Clk_period;
		Addr <=  "0011010000110";
		Trees_din <= x"ffeb1b85";
		wait for Clk_period;
		Addr <=  "0011010000111";
		Trees_din <= x"008b1b85";
		wait for Clk_period;
		Addr <=  "0011010001000";
		Trees_din <= x"1400e304";
		wait for Clk_period;
		Addr <=  "0011010001001";
		Trees_din <= x"00151b85";
		wait for Clk_period;
		Addr <=  "0011010001010";
		Trees_din <= x"ff131b85";
		wait for Clk_period;
		Addr <=  "0011010001011";
		Trees_din <= x"08003b08";
		wait for Clk_period;
		Addr <=  "0011010001100";
		Trees_din <= x"09010a04";
		wait for Clk_period;
		Addr <=  "0011010001101";
		Trees_din <= x"00b81b85";
		wait for Clk_period;
		Addr <=  "0011010001110";
		Trees_din <= x"ffad1b85";
		wait for Clk_period;
		Addr <=  "0011010001111";
		Trees_din <= x"19000004";
		wait for Clk_period;
		Addr <=  "0011010010000";
		Trees_din <= x"ff9e1b85";
		wait for Clk_period;
		Addr <=  "0011010010001";
		Trees_din <= x"001c1b85";
		wait for Clk_period;
		Addr <=  "0011010010010";
		Trees_din <= x"0209d010";
		wait for Clk_period;
		Addr <=  "0011010010011";
		Trees_din <= x"19000108";
		wait for Clk_period;
		Addr <=  "0011010010100";
		Trees_din <= x"0c009904";
		wait for Clk_period;
		Addr <=  "0011010010101";
		Trees_din <= x"001b1b85";
		wait for Clk_period;
		Addr <=  "0011010010110";
		Trees_din <= x"00b31b85";
		wait for Clk_period;
		Addr <=  "0011010010111";
		Trees_din <= x"06ff7604";
		wait for Clk_period;
		Addr <=  "0011010011000";
		Trees_din <= x"ffc81b85";
		wait for Clk_period;
		Addr <=  "0011010011001";
		Trees_din <= x"00941b85";
		wait for Clk_period;
		Addr <=  "0011010011010";
		Trees_din <= x"0e003104";
		wait for Clk_period;
		Addr <=  "0011010011011";
		Trees_din <= x"ff601b85";
		wait for Clk_period;
		Addr <=  "0011010011100";
		Trees_din <= x"ffff1b85";
		wait for Clk_period;
		Addr <=  "0011010011101";
		Trees_din <= x"04054320";
		wait for Clk_period;
		Addr <=  "0011010011110";
		Trees_din <= x"02046810";
		wait for Clk_period;
		Addr <=  "0011010011111";
		Trees_din <= x"010ab108";
		wait for Clk_period;
		Addr <=  "0011010100000";
		Trees_din <= x"10004104";
		wait for Clk_period;
		Addr <=  "0011010100001";
		Trees_din <= x"00421b85";
		wait for Clk_period;
		Addr <=  "0011010100010";
		Trees_din <= x"ffcc1b85";
		wait for Clk_period;
		Addr <=  "0011010100011";
		Trees_din <= x"05f5e804";
		wait for Clk_period;
		Addr <=  "0011010100100";
		Trees_din <= x"00081b85";
		wait for Clk_period;
		Addr <=  "0011010100101";
		Trees_din <= x"00601b85";
		wait for Clk_period;
		Addr <=  "0011010100110";
		Trees_din <= x"06019008";
		wait for Clk_period;
		Addr <=  "0011010100111";
		Trees_din <= x"04020704";
		wait for Clk_period;
		Addr <=  "0011010101000";
		Trees_din <= x"ffd31b85";
		wait for Clk_period;
		Addr <=  "0011010101001";
		Trees_din <= x"00471b85";
		wait for Clk_period;
		Addr <=  "0011010101010";
		Trees_din <= x"0d000204";
		wait for Clk_period;
		Addr <=  "0011010101011";
		Trees_din <= x"ff871b85";
		wait for Clk_period;
		Addr <=  "0011010101100";
		Trees_din <= x"00341b85";
		wait for Clk_period;
		Addr <=  "0011010101101";
		Trees_din <= x"1500450c";
		wait for Clk_period;
		Addr <=  "0011010101110";
		Trees_din <= x"19000008";
		wait for Clk_period;
		Addr <=  "0011010101111";
		Trees_din <= x"12007404";
		wait for Clk_period;
		Addr <=  "0011010110000";
		Trees_din <= x"00ea1b85";
		wait for Clk_period;
		Addr <=  "0011010110001";
		Trees_din <= x"00421b85";
		wait for Clk_period;
		Addr <=  "0011010110010";
		Trees_din <= x"ffff1b85";
		wait for Clk_period;
		Addr <=  "0011010110011";
		Trees_din <= x"ffd51b85";
		wait for Clk_period;
		Addr <=  "0011010110100";
		Trees_din <= x"1403fe40";
		wait for Clk_period;
		Addr <=  "0011010110101";
		Trees_din <= x"04fdb120";
		wait for Clk_period;
		Addr <=  "0011010110110";
		Trees_din <= x"0e002f10";
		wait for Clk_period;
		Addr <=  "0011010110111";
		Trees_din <= x"1802b308";
		wait for Clk_period;
		Addr <=  "0011010111000";
		Trees_din <= x"15003004";
		wait for Clk_period;
		Addr <=  "0011010111001";
		Trees_din <= x"ff921b85";
		wait for Clk_period;
		Addr <=  "0011010111010";
		Trees_din <= x"00231b85";
		wait for Clk_period;
		Addr <=  "0011010111011";
		Trees_din <= x"1101f304";
		wait for Clk_period;
		Addr <=  "0011010111100";
		Trees_din <= x"00b81b85";
		wait for Clk_period;
		Addr <=  "0011010111101";
		Trees_din <= x"000a1b85";
		wait for Clk_period;
		Addr <=  "0011010111110";
		Trees_din <= x"0703ea08";
		wait for Clk_period;
		Addr <=  "0011010111111";
		Trees_din <= x"01114c04";
		wait for Clk_period;
		Addr <=  "0011011000000";
		Trees_din <= x"ff8d1b85";
		wait for Clk_period;
		Addr <=  "0011011000001";
		Trees_din <= x"00691b85";
		wait for Clk_period;
		Addr <=  "0011011000010";
		Trees_din <= x"13019c04";
		wait for Clk_period;
		Addr <=  "0011011000011";
		Trees_din <= x"007d1b85";
		wait for Clk_period;
		Addr <=  "0011011000100";
		Trees_din <= x"fff21b85";
		wait for Clk_period;
		Addr <=  "0011011000101";
		Trees_din <= x"04ffdd10";
		wait for Clk_period;
		Addr <=  "0011011000110";
		Trees_din <= x"0d020508";
		wait for Clk_period;
		Addr <=  "0011011000111";
		Trees_din <= x"02076e04";
		wait for Clk_period;
		Addr <=  "0011011001000";
		Trees_din <= x"00291b85";
		wait for Clk_period;
		Addr <=  "0011011001001";
		Trees_din <= x"00ac1b85";
		wait for Clk_period;
		Addr <=  "0011011001010";
		Trees_din <= x"09008a04";
		wait for Clk_period;
		Addr <=  "0011011001011";
		Trees_din <= x"006e1b85";
		wait for Clk_period;
		Addr <=  "0011011001100";
		Trees_din <= x"ffc41b85";
		wait for Clk_period;
		Addr <=  "0011011001101";
		Trees_din <= x"0b007e08";
		wait for Clk_period;
		Addr <=  "0011011001110";
		Trees_din <= x"12007d04";
		wait for Clk_period;
		Addr <=  "0011011001111";
		Trees_din <= x"ffe01b85";
		wait for Clk_period;
		Addr <=  "0011011010000";
		Trees_din <= x"00841b85";
		wait for Clk_period;
		Addr <=  "0011011010001";
		Trees_din <= x"05f52b04";
		wait for Clk_period;
		Addr <=  "0011011010010";
		Trees_din <= x"ffdd1b85";
		wait for Clk_period;
		Addr <=  "0011011010011";
		Trees_din <= x"ff461b85";
		wait for Clk_period;
		Addr <=  "0011011010100";
		Trees_din <= x"0800440c";
		wait for Clk_period;
		Addr <=  "0011011010101";
		Trees_din <= x"02056b04";
		wait for Clk_period;
		Addr <=  "0011011010110";
		Trees_din <= x"ffee1b85";
		wait for Clk_period;
		Addr <=  "0011011010111";
		Trees_din <= x"15003a04";
		wait for Clk_period;
		Addr <=  "0011011011000";
		Trees_din <= x"ffcd1b85";
		wait for Clk_period;
		Addr <=  "0011011011001";
		Trees_din <= x"ff101b85";
		wait for Clk_period;
		Addr <=  "0011011011010";
		Trees_din <= x"1403ff04";
		wait for Clk_period;
		Addr <=  "0011011011011";
		Trees_din <= x"ff621b85";
		wait for Clk_period;
		Addr <=  "0011011011100";
		Trees_din <= x"1403ff04";
		wait for Clk_period;
		Addr <=  "0011011011101";
		Trees_din <= x"00a71b85";
		wait for Clk_period;
		Addr <=  "0011011011110";
		Trees_din <= x"0b006b04";
		wait for Clk_period;
		Addr <=  "0011011011111";
		Trees_din <= x"ffa41b85";
		wait for Clk_period;
		Addr <=  "0011011100000";
		Trees_din <= x"00321b85";
		wait for Clk_period;
		Addr <=  "0011011100001";
		Trees_din <= x"0111f868";
		wait for Clk_period;
		Addr <=  "0011011100010";
		Trees_din <= x"1402372c";
		wait for Clk_period;
		Addr <=  "0011011100011";
		Trees_din <= x"08002d0c";
		wait for Clk_period;
		Addr <=  "0011011100100";
		Trees_din <= x"05f3ca04";
		wait for Clk_period;
		Addr <=  "0011011100101";
		Trees_din <= x"002b1ca1";
		wait for Clk_period;
		Addr <=  "0011011100110";
		Trees_din <= x"12007e04";
		wait for Clk_period;
		Addr <=  "0011011100111";
		Trees_din <= x"ffdb1ca1";
		wait for Clk_period;
		Addr <=  "0011011101000";
		Trees_din <= x"ff661ca1";
		wait for Clk_period;
		Addr <=  "0011011101001";
		Trees_din <= x"19000b10";
		wait for Clk_period;
		Addr <=  "0011011101010";
		Trees_din <= x"1f028608";
		wait for Clk_period;
		Addr <=  "0011011101011";
		Trees_din <= x"1c028204";
		wait for Clk_period;
		Addr <=  "0011011101100";
		Trees_din <= x"00051ca1";
		wait for Clk_period;
		Addr <=  "0011011101101";
		Trees_din <= x"009d1ca1";
		wait for Clk_period;
		Addr <=  "0011011101110";
		Trees_din <= x"19000004";
		wait for Clk_period;
		Addr <=  "0011011101111";
		Trees_din <= x"002a1ca1";
		wait for Clk_period;
		Addr <=  "0011011110000";
		Trees_din <= x"ff771ca1";
		wait for Clk_period;
		Addr <=  "0011011110001";
		Trees_din <= x"1a018708";
		wait for Clk_period;
		Addr <=  "0011011110010";
		Trees_din <= x"03fa8604";
		wait for Clk_period;
		Addr <=  "0011011110011";
		Trees_din <= x"00cc1ca1";
		wait for Clk_period;
		Addr <=  "0011011110100";
		Trees_din <= x"00201ca1";
		wait for Clk_period;
		Addr <=  "0011011110101";
		Trees_din <= x"010acf04";
		wait for Clk_period;
		Addr <=  "0011011110110";
		Trees_din <= x"ffa41ca1";
		wait for Clk_period;
		Addr <=  "0011011110111";
		Trees_din <= x"004a1ca1";
		wait for Clk_period;
		Addr <=  "0011011111000";
		Trees_din <= x"18006b20";
		wait for Clk_period;
		Addr <=  "0011011111001";
		Trees_din <= x"1b027410";
		wait for Clk_period;
		Addr <=  "0011011111010";
		Trees_din <= x"0405f108";
		wait for Clk_period;
		Addr <=  "0011011111011";
		Trees_din <= x"05f56304";
		wait for Clk_period;
		Addr <=  "0011011111100";
		Trees_din <= x"00161ca1";
		wait for Clk_period;
		Addr <=  "0011011111101";
		Trees_din <= x"ffed1ca1";
		wait for Clk_period;
		Addr <=  "0011011111110";
		Trees_din <= x"0a004604";
		wait for Clk_period;
		Addr <=  "0011011111111";
		Trees_din <= x"00ab1ca1";
		wait for Clk_period;
		Addr <=  "0011100000000";
		Trees_din <= x"00071ca1";
		wait for Clk_period;
		Addr <=  "0011100000001";
		Trees_din <= x"07fa1c08";
		wait for Clk_period;
		Addr <=  "0011100000010";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0011100000011";
		Trees_din <= x"fffa1ca1";
		wait for Clk_period;
		Addr <=  "0011100000100";
		Trees_din <= x"00c91ca1";
		wait for Clk_period;
		Addr <=  "0011100000101";
		Trees_din <= x"17f83204";
		wait for Clk_period;
		Addr <=  "0011100000110";
		Trees_din <= x"006b1ca1";
		wait for Clk_period;
		Addr <=  "0011100000111";
		Trees_din <= x"ffe81ca1";
		wait for Clk_period;
		Addr <=  "0011100001000";
		Trees_din <= x"1403f810";
		wait for Clk_period;
		Addr <=  "0011100001001";
		Trees_din <= x"03f86708";
		wait for Clk_period;
		Addr <=  "0011100001010";
		Trees_din <= x"16007004";
		wait for Clk_period;
		Addr <=  "0011100001011";
		Trees_din <= x"fff71ca1";
		wait for Clk_period;
		Addr <=  "0011100001100";
		Trees_din <= x"ffb41ca1";
		wait for Clk_period;
		Addr <=  "0011100001101";
		Trees_din <= x"0f008604";
		wait for Clk_period;
		Addr <=  "0011100001110";
		Trees_din <= x"00241ca1";
		wait for Clk_period;
		Addr <=  "0011100001111";
		Trees_din <= x"ffd71ca1";
		wait for Clk_period;
		Addr <=  "0011100010000";
		Trees_din <= x"0d018e08";
		wait for Clk_period;
		Addr <=  "0011100010001";
		Trees_din <= x"1100dd04";
		wait for Clk_period;
		Addr <=  "0011100010010";
		Trees_din <= x"001a1ca1";
		wait for Clk_period;
		Addr <=  "0011100010011";
		Trees_din <= x"ff6b1ca1";
		wait for Clk_period;
		Addr <=  "0011100010100";
		Trees_din <= x"00691ca1";
		wait for Clk_period;
		Addr <=  "0011100010101";
		Trees_din <= x"000e1910";
		wait for Clk_period;
		Addr <=  "0011100010110";
		Trees_din <= x"08003008";
		wait for Clk_period;
		Addr <=  "0011100010111";
		Trees_din <= x"0c00af04";
		wait for Clk_period;
		Addr <=  "0011100011000";
		Trees_din <= x"00591ca1";
		wait for Clk_period;
		Addr <=  "0011100011001";
		Trees_din <= x"ffbd1ca1";
		wait for Clk_period;
		Addr <=  "0011100011010";
		Trees_din <= x"16009104";
		wait for Clk_period;
		Addr <=  "0011100011011";
		Trees_din <= x"008d1ca1";
		wait for Clk_period;
		Addr <=  "0011100011100";
		Trees_din <= x"00241ca1";
		wait for Clk_period;
		Addr <=  "0011100011101";
		Trees_din <= x"08003f0c";
		wait for Clk_period;
		Addr <=  "0011100011110";
		Trees_din <= x"08003704";
		wait for Clk_period;
		Addr <=  "0011100011111";
		Trees_din <= x"00551ca1";
		wait for Clk_period;
		Addr <=  "0011100100000";
		Trees_din <= x"17f7b504";
		wait for Clk_period;
		Addr <=  "0011100100001";
		Trees_din <= x"ff801ca1";
		wait for Clk_period;
		Addr <=  "0011100100010";
		Trees_din <= x"00071ca1";
		wait for Clk_period;
		Addr <=  "0011100100011";
		Trees_din <= x"0f008d08";
		wait for Clk_period;
		Addr <=  "0011100100100";
		Trees_din <= x"18000904";
		wait for Clk_period;
		Addr <=  "0011100100101";
		Trees_din <= x"ffde1ca1";
		wait for Clk_period;
		Addr <=  "0011100100110";
		Trees_din <= x"00741ca1";
		wait for Clk_period;
		Addr <=  "0011100100111";
		Trees_din <= x"ffcf1ca1";
		wait for Clk_period;
		Addr <=  "0011100101000";
		Trees_din <= x"0106bc38";
		wait for Clk_period;
		Addr <=  "0011100101001";
		Trees_din <= x"19000124";
		wait for Clk_period;
		Addr <=  "0011100101010";
		Trees_din <= x"16008220";
		wait for Clk_period;
		Addr <=  "0011100101011";
		Trees_din <= x"12007310";
		wait for Clk_period;
		Addr <=  "0011100101100";
		Trees_din <= x"0105ce08";
		wait for Clk_period;
		Addr <=  "0011100101101";
		Trees_din <= x"16006904";
		wait for Clk_period;
		Addr <=  "0011100101110";
		Trees_din <= x"00981df5";
		wait for Clk_period;
		Addr <=  "0011100101111";
		Trees_din <= x"ffc81df5";
		wait for Clk_period;
		Addr <=  "0011100110000";
		Trees_din <= x"1100d204";
		wait for Clk_period;
		Addr <=  "0011100110001";
		Trees_din <= x"00511df5";
		wait for Clk_period;
		Addr <=  "0011100110010";
		Trees_din <= x"00fc1df5";
		wait for Clk_period;
		Addr <=  "0011100110011";
		Trees_din <= x"0c00b308";
		wait for Clk_period;
		Addr <=  "0011100110100";
		Trees_din <= x"07040e04";
		wait for Clk_period;
		Addr <=  "0011100110101";
		Trees_din <= x"ff6f1df5";
		wait for Clk_period;
		Addr <=  "0011100110110";
		Trees_din <= x"00021df5";
		wait for Clk_period;
		Addr <=  "0011100110111";
		Trees_din <= x"11017c04";
		wait for Clk_period;
		Addr <=  "0011100111000";
		Trees_din <= x"00531df5";
		wait for Clk_period;
		Addr <=  "0011100111001";
		Trees_din <= x"ff881df5";
		wait for Clk_period;
		Addr <=  "0011100111010";
		Trees_din <= x"ff7c1df5";
		wait for Clk_period;
		Addr <=  "0011100111011";
		Trees_din <= x"0d02050c";
		wait for Clk_period;
		Addr <=  "0011100111100";
		Trees_din <= x"05fd0304";
		wait for Clk_period;
		Addr <=  "0011100111101";
		Trees_din <= x"ff631df5";
		wait for Clk_period;
		Addr <=  "0011100111110";
		Trees_din <= x"0600c004";
		wait for Clk_period;
		Addr <=  "0011100111111";
		Trees_din <= x"00301df5";
		wait for Clk_period;
		Addr <=  "0011101000000";
		Trees_din <= x"ff9f1df5";
		wait for Clk_period;
		Addr <=  "0011101000001";
		Trees_din <= x"1af9f404";
		wait for Clk_period;
		Addr <=  "0011101000010";
		Trees_din <= x"007b1df5";
		wait for Clk_period;
		Addr <=  "0011101000011";
		Trees_din <= x"00011df5";
		wait for Clk_period;
		Addr <=  "0011101000100";
		Trees_din <= x"0601ac40";
		wait for Clk_period;
		Addr <=  "0011101000101";
		Trees_din <= x"0a005220";
		wait for Clk_period;
		Addr <=  "0011101000110";
		Trees_din <= x"17f74210";
		wait for Clk_period;
		Addr <=  "0011101000111";
		Trees_din <= x"0900ef08";
		wait for Clk_period;
		Addr <=  "0011101001000";
		Trees_din <= x"0e002e04";
		wait for Clk_period;
		Addr <=  "0011101001001";
		Trees_din <= x"ff831df5";
		wait for Clk_period;
		Addr <=  "0011101001010";
		Trees_din <= x"ffe71df5";
		wait for Clk_period;
		Addr <=  "0011101001011";
		Trees_din <= x"02046804";
		wait for Clk_period;
		Addr <=  "0011101001100";
		Trees_din <= x"009d1df5";
		wait for Clk_period;
		Addr <=  "0011101001101";
		Trees_din <= x"00001df5";
		wait for Clk_period;
		Addr <=  "0011101001110";
		Trees_din <= x"1b025908";
		wait for Clk_period;
		Addr <=  "0011101001111";
		Trees_din <= x"0e003e04";
		wait for Clk_period;
		Addr <=  "0011101010000";
		Trees_din <= x"005c1df5";
		wait for Clk_period;
		Addr <=  "0011101010001";
		Trees_din <= x"ffd91df5";
		wait for Clk_period;
		Addr <=  "0011101010010";
		Trees_din <= x"03f86704";
		wait for Clk_period;
		Addr <=  "0011101010011";
		Trees_din <= x"ffeb1df5";
		wait for Clk_period;
		Addr <=  "0011101010100";
		Trees_din <= x"00101df5";
		wait for Clk_period;
		Addr <=  "0011101010101";
		Trees_din <= x"04ffbc10";
		wait for Clk_period;
		Addr <=  "0011101010110";
		Trees_din <= x"07fb7208";
		wait for Clk_period;
		Addr <=  "0011101010111";
		Trees_din <= x"07f99f04";
		wait for Clk_period;
		Addr <=  "0011101011000";
		Trees_din <= x"002c1df5";
		wait for Clk_period;
		Addr <=  "0011101011001";
		Trees_din <= x"ff5b1df5";
		wait for Clk_period;
		Addr <=  "0011101011010";
		Trees_din <= x"1e027f04";
		wait for Clk_period;
		Addr <=  "0011101011011";
		Trees_din <= x"006c1df5";
		wait for Clk_period;
		Addr <=  "0011101011100";
		Trees_din <= x"ffe51df5";
		wait for Clk_period;
		Addr <=  "0011101011101";
		Trees_din <= x"07f77b08";
		wait for Clk_period;
		Addr <=  "0011101011110";
		Trees_din <= x"1403f604";
		wait for Clk_period;
		Addr <=  "0011101011111";
		Trees_din <= x"ff961df5";
		wait for Clk_period;
		Addr <=  "0011101100000";
		Trees_din <= x"002e1df5";
		wait for Clk_period;
		Addr <=  "0011101100001";
		Trees_din <= x"05f25604";
		wait for Clk_period;
		Addr <=  "0011101100010";
		Trees_din <= x"ffd11df5";
		wait for Clk_period;
		Addr <=  "0011101100011";
		Trees_din <= x"00a01df5";
		wait for Clk_period;
		Addr <=  "0011101100100";
		Trees_din <= x"0a005020";
		wait for Clk_period;
		Addr <=  "0011101100101";
		Trees_din <= x"0c00c810";
		wait for Clk_period;
		Addr <=  "0011101100110";
		Trees_din <= x"12007c08";
		wait for Clk_period;
		Addr <=  "0011101100111";
		Trees_din <= x"1d025c04";
		wait for Clk_period;
		Addr <=  "0011101101000";
		Trees_din <= x"00661df5";
		wait for Clk_period;
		Addr <=  "0011101101001";
		Trees_din <= x"ffff1df5";
		wait for Clk_period;
		Addr <=  "0011101101010";
		Trees_din <= x"0f000304";
		wait for Clk_period;
		Addr <=  "0011101101011";
		Trees_din <= x"ffe91df5";
		wait for Clk_period;
		Addr <=  "0011101101100";
		Trees_din <= x"00c71df5";
		wait for Clk_period;
		Addr <=  "0011101101101";
		Trees_din <= x"0c00ec08";
		wait for Clk_period;
		Addr <=  "0011101101110";
		Trees_din <= x"1b026904";
		wait for Clk_period;
		Addr <=  "0011101101111";
		Trees_din <= x"00311df5";
		wait for Clk_period;
		Addr <=  "0011101110000";
		Trees_din <= x"ff801df5";
		wait for Clk_period;
		Addr <=  "0011101110001";
		Trees_din <= x"07fb8104";
		wait for Clk_period;
		Addr <=  "0011101110010";
		Trees_din <= x"00af1df5";
		wait for Clk_period;
		Addr <=  "0011101110011";
		Trees_din <= x"ffdc1df5";
		wait for Clk_period;
		Addr <=  "0011101110100";
		Trees_din <= x"12007d08";
		wait for Clk_period;
		Addr <=  "0011101110101";
		Trees_din <= x"0f000104";
		wait for Clk_period;
		Addr <=  "0011101110110";
		Trees_din <= x"00781df5";
		wait for Clk_period;
		Addr <=  "0011101110111";
		Trees_din <= x"ffcf1df5";
		wait for Clk_period;
		Addr <=  "0011101111000";
		Trees_din <= x"1403b704";
		wait for Clk_period;
		Addr <=  "0011101111001";
		Trees_din <= x"002d1df5";
		wait for Clk_period;
		Addr <=  "0011101111010";
		Trees_din <= x"06044604";
		wait for Clk_period;
		Addr <=  "0011101111011";
		Trees_din <= x"ff351df5";
		wait for Clk_period;
		Addr <=  "0011101111100";
		Trees_din <= x"00241df5";
		wait for Clk_period;
		Addr <=  "0011101111101";
		Trees_din <= x"0111f840";
		wait for Clk_period;
		Addr <=  "0011101111110";
		Trees_din <= x"01ffc904";
		wait for Clk_period;
		Addr <=  "0011101111111";
		Trees_din <= x"ff881ec9";
		wait for Clk_period;
		Addr <=  "0011110000000";
		Trees_din <= x"03f47620";
		wait for Clk_period;
		Addr <=  "0011110000001";
		Trees_din <= x"0900e310";
		wait for Clk_period;
		Addr <=  "0011110000010";
		Trees_din <= x"0b008608";
		wait for Clk_period;
		Addr <=  "0011110000011";
		Trees_din <= x"19000304";
		wait for Clk_period;
		Addr <=  "0011110000100";
		Trees_din <= x"00a61ec9";
		wait for Clk_period;
		Addr <=  "0011110000101";
		Trees_din <= x"00111ec9";
		wait for Clk_period;
		Addr <=  "0011110000110";
		Trees_din <= x"12009904";
		wait for Clk_period;
		Addr <=  "0011110000111";
		Trees_din <= x"ff8a1ec9";
		wait for Clk_period;
		Addr <=  "0011110001000";
		Trees_din <= x"00501ec9";
		wait for Clk_period;
		Addr <=  "0011110001001";
		Trees_din <= x"0e002408";
		wait for Clk_period;
		Addr <=  "0011110001010";
		Trees_din <= x"1c024704";
		wait for Clk_period;
		Addr <=  "0011110001011";
		Trees_din <= x"00a31ec9";
		wait for Clk_period;
		Addr <=  "0011110001100";
		Trees_din <= x"ffcb1ec9";
		wait for Clk_period;
		Addr <=  "0011110001101";
		Trees_din <= x"1afb2804";
		wait for Clk_period;
		Addr <=  "0011110001110";
		Trees_din <= x"002d1ec9";
		wait for Clk_period;
		Addr <=  "0011110001111";
		Trees_din <= x"ff761ec9";
		wait for Clk_period;
		Addr <=  "0011110010000";
		Trees_din <= x"04020710";
		wait for Clk_period;
		Addr <=  "0011110010001";
		Trees_din <= x"020ba008";
		wait for Clk_period;
		Addr <=  "0011110010010";
		Trees_din <= x"03f49404";
		wait for Clk_period;
		Addr <=  "0011110010011";
		Trees_din <= x"ff581ec9";
		wait for Clk_period;
		Addr <=  "0011110010100";
		Trees_din <= x"fffb1ec9";
		wait for Clk_period;
		Addr <=  "0011110010101";
		Trees_din <= x"04009f04";
		wait for Clk_period;
		Addr <=  "0011110010110";
		Trees_din <= x"00b01ec9";
		wait for Clk_period;
		Addr <=  "0011110010111";
		Trees_din <= x"ffaa1ec9";
		wait for Clk_period;
		Addr <=  "0011110011000";
		Trees_din <= x"1c028508";
		wait for Clk_period;
		Addr <=  "0011110011001";
		Trees_din <= x"06024704";
		wait for Clk_period;
		Addr <=  "0011110011010";
		Trees_din <= x"00421ec9";
		wait for Clk_period;
		Addr <=  "0011110011011";
		Trees_din <= x"ffd51ec9";
		wait for Clk_period;
		Addr <=  "0011110011100";
		Trees_din <= x"ff6c1ec9";
		wait for Clk_period;
		Addr <=  "0011110011101";
		Trees_din <= x"07f87a1c";
		wait for Clk_period;
		Addr <=  "0011110011110";
		Trees_din <= x"05f2c114";
		wait for Clk_period;
		Addr <=  "0011110011111";
		Trees_din <= x"07f70a0c";
		wait for Clk_period;
		Addr <=  "0011110100000";
		Trees_din <= x"08003f08";
		wait for Clk_period;
		Addr <=  "0011110100001";
		Trees_din <= x"10004904";
		wait for Clk_period;
		Addr <=  "0011110100010";
		Trees_din <= x"ffcf1ec9";
		wait for Clk_period;
		Addr <=  "0011110100011";
		Trees_din <= x"fff71ec9";
		wait for Clk_period;
		Addr <=  "0011110100100";
		Trees_din <= x"00611ec9";
		wait for Clk_period;
		Addr <=  "0011110100101";
		Trees_din <= x"0c00a404";
		wait for Clk_period;
		Addr <=  "0011110100110";
		Trees_din <= x"00011ec9";
		wait for Clk_period;
		Addr <=  "0011110100111";
		Trees_din <= x"ff7a1ec9";
		wait for Clk_period;
		Addr <=  "0011110101000";
		Trees_din <= x"0400c804";
		wait for Clk_period;
		Addr <=  "0011110101001";
		Trees_din <= x"006a1ec9";
		wait for Clk_period;
		Addr <=  "0011110101010";
		Trees_din <= x"00091ec9";
		wait for Clk_period;
		Addr <=  "0011110101011";
		Trees_din <= x"06fbe10c";
		wait for Clk_period;
		Addr <=  "0011110101100";
		Trees_din <= x"06fb7508";
		wait for Clk_period;
		Addr <=  "0011110101101";
		Trees_din <= x"08004404";
		wait for Clk_period;
		Addr <=  "0011110101110";
		Trees_din <= x"00671ec9";
		wait for Clk_period;
		Addr <=  "0011110101111";
		Trees_din <= x"00161ec9";
		wait for Clk_period;
		Addr <=  "0011110110000";
		Trees_din <= x"ffbc1ec9";
		wait for Clk_period;
		Addr <=  "0011110110001";
		Trees_din <= x"008b1ec9";
		wait for Clk_period;
		Addr <=  "0011110110010";
		Trees_din <= x"0111f844";
		wait for Clk_period;
		Addr <=  "0011110110011";
		Trees_din <= x"1dfd6220";
		wait for Clk_period;
		Addr <=  "0011110110100";
		Trees_din <= x"03f9bb14";
		wait for Clk_period;
		Addr <=  "0011110110101";
		Trees_din <= x"15003d0c";
		wait for Clk_period;
		Addr <=  "0011110110110";
		Trees_din <= x"14029004";
		wait for Clk_period;
		Addr <=  "0011110110111";
		Trees_din <= x"00b51f9d";
		wait for Clk_period;
		Addr <=  "0011110111000";
		Trees_din <= x"0a003e04";
		wait for Clk_period;
		Addr <=  "0011110111001";
		Trees_din <= x"00781f9d";
		wait for Clk_period;
		Addr <=  "0011110111010";
		Trees_din <= x"ffc51f9d";
		wait for Clk_period;
		Addr <=  "0011110111011";
		Trees_din <= x"12007004";
		wait for Clk_period;
		Addr <=  "0011110111100";
		Trees_din <= x"00231f9d";
		wait for Clk_period;
		Addr <=  "0011110111101";
		Trees_din <= x"ff9d1f9d";
		wait for Clk_period;
		Addr <=  "0011110111110";
		Trees_din <= x"1ff9b004";
		wait for Clk_period;
		Addr <=  "0011110111111";
		Trees_din <= x"004a1f9d";
		wait for Clk_period;
		Addr <=  "0011111000000";
		Trees_din <= x"03fb8604";
		wait for Clk_period;
		Addr <=  "0011111000001";
		Trees_din <= x"ff7f1f9d";
		wait for Clk_period;
		Addr <=  "0011111000010";
		Trees_din <= x"fff91f9d";
		wait for Clk_period;
		Addr <=  "0011111000011";
		Trees_din <= x"1dfdb404";
		wait for Clk_period;
		Addr <=  "0011111000100";
		Trees_din <= x"ff7d1f9d";
		wait for Clk_period;
		Addr <=  "0011111000101";
		Trees_din <= x"0c00f410";
		wait for Clk_period;
		Addr <=  "0011111000110";
		Trees_din <= x"0c00cb08";
		wait for Clk_period;
		Addr <=  "0011111000111";
		Trees_din <= x"15003504";
		wait for Clk_period;
		Addr <=  "0011111001000";
		Trees_din <= x"00341f9d";
		wait for Clk_period;
		Addr <=  "0011111001001";
		Trees_din <= x"fffe1f9d";
		wait for Clk_period;
		Addr <=  "0011111001010";
		Trees_din <= x"0b009d04";
		wait for Clk_period;
		Addr <=  "0011111001011";
		Trees_din <= x"ffcc1f9d";
		wait for Clk_period;
		Addr <=  "0011111001100";
		Trees_din <= x"003b1f9d";
		wait for Clk_period;
		Addr <=  "0011111001101";
		Trees_din <= x"10002f08";
		wait for Clk_period;
		Addr <=  "0011111001110";
		Trees_din <= x"05f46b04";
		wait for Clk_period;
		Addr <=  "0011111001111";
		Trees_din <= x"005c1f9d";
		wait for Clk_period;
		Addr <=  "0011111010000";
		Trees_din <= x"ffa81f9d";
		wait for Clk_period;
		Addr <=  "0011111010001";
		Trees_din <= x"000dd104";
		wait for Clk_period;
		Addr <=  "0011111010010";
		Trees_din <= x"008e1f9d";
		wait for Clk_period;
		Addr <=  "0011111010011";
		Trees_din <= x"ffa61f9d";
		wait for Clk_period;
		Addr <=  "0011111010100";
		Trees_din <= x"07f87a18";
		wait for Clk_period;
		Addr <=  "0011111010101";
		Trees_din <= x"05f2c110";
		wait for Clk_period;
		Addr <=  "0011111010110";
		Trees_din <= x"07f70a08";
		wait for Clk_period;
		Addr <=  "0011111010111";
		Trees_din <= x"08003f04";
		wait for Clk_period;
		Addr <=  "0011111011000";
		Trees_din <= x"ffdc1f9d";
		wait for Clk_period;
		Addr <=  "0011111011001";
		Trees_din <= x"005c1f9d";
		wait for Clk_period;
		Addr <=  "0011111011010";
		Trees_din <= x"0c00a404";
		wait for Clk_period;
		Addr <=  "0011111011011";
		Trees_din <= x"00011f9d";
		wait for Clk_period;
		Addr <=  "0011111011100";
		Trees_din <= x"ff871f9d";
		wait for Clk_period;
		Addr <=  "0011111011101";
		Trees_din <= x"0e003904";
		wait for Clk_period;
		Addr <=  "0011111011110";
		Trees_din <= x"00661f9d";
		wait for Clk_period;
		Addr <=  "0011111011111";
		Trees_din <= x"00081f9d";
		wait for Clk_period;
		Addr <=  "0011111100000";
		Trees_din <= x"06fbe10c";
		wait for Clk_period;
		Addr <=  "0011111100001";
		Trees_din <= x"06fb7508";
		wait for Clk_period;
		Addr <=  "0011111100010";
		Trees_din <= x"08004404";
		wait for Clk_period;
		Addr <=  "0011111100011";
		Trees_din <= x"00631f9d";
		wait for Clk_period;
		Addr <=  "0011111100100";
		Trees_din <= x"00151f9d";
		wait for Clk_period;
		Addr <=  "0011111100101";
		Trees_din <= x"ffc21f9d";
		wait for Clk_period;
		Addr <=  "0011111100110";
		Trees_din <= x"00881f9d";
		wait for Clk_period;
		Addr <=  "0011111100111";
		Trees_din <= x"16009160";
		wait for Clk_period;
		Addr <=  "0011111101000";
		Trees_din <= x"0c007b24";
		wait for Clk_period;
		Addr <=  "0011111101001";
		Trees_din <= x"000c1218";
		wait for Clk_period;
		Addr <=  "0011111101010";
		Trees_din <= x"1500410c";
		wait for Clk_period;
		Addr <=  "0011111101011";
		Trees_din <= x"010b8304";
		wait for Clk_period;
		Addr <=  "0011111101100";
		Trees_din <= x"ff8e20d1";
		wait for Clk_period;
		Addr <=  "0011111101101";
		Trees_din <= x"05f48f04";
		wait for Clk_period;
		Addr <=  "0011111101110";
		Trees_din <= x"ffd820d1";
		wait for Clk_period;
		Addr <=  "0011111101111";
		Trees_din <= x"006720d1";
		wait for Clk_period;
		Addr <=  "0011111110000";
		Trees_din <= x"05f46b04";
		wait for Clk_period;
		Addr <=  "0011111110001";
		Trees_din <= x"002b20d1";
		wait for Clk_period;
		Addr <=  "0011111110010";
		Trees_din <= x"17f7b504";
		wait for Clk_period;
		Addr <=  "0011111110011";
		Trees_din <= x"ff2320d1";
		wait for Clk_period;
		Addr <=  "0011111110100";
		Trees_din <= x"ffba20d1";
		wait for Clk_period;
		Addr <=  "0011111110101";
		Trees_din <= x"03f66004";
		wait for Clk_period;
		Addr <=  "0011111110110";
		Trees_din <= x"ff9e20d1";
		wait for Clk_period;
		Addr <=  "0011111110111";
		Trees_din <= x"000de204";
		wait for Clk_period;
		Addr <=  "0011111111000";
		Trees_din <= x"009120d1";
		wait for Clk_period;
		Addr <=  "0011111111001";
		Trees_din <= x"002120d1";
		wait for Clk_period;
		Addr <=  "0011111111010";
		Trees_din <= x"11018520";
		wait for Clk_period;
		Addr <=  "0011111111011";
		Trees_din <= x"21000010";
		wait for Clk_period;
		Addr <=  "0011111111100";
		Trees_din <= x"0d000308";
		wait for Clk_period;
		Addr <=  "0011111111101";
		Trees_din <= x"0e003804";
		wait for Clk_period;
		Addr <=  "0011111111110";
		Trees_din <= x"006920d1";
		wait for Clk_period;
		Addr <=  "0011111111111";
		Trees_din <= x"ffc320d1";
		wait for Clk_period;
		Addr <=  "0100000000000";
		Trees_din <= x"14021504";
		wait for Clk_period;
		Addr <=  "0100000000001";
		Trees_din <= x"005620d1";
		wait for Clk_period;
		Addr <=  "0100000000010";
		Trees_din <= x"000b20d1";
		wait for Clk_period;
		Addr <=  "0100000000011";
		Trees_din <= x"04fdc308";
		wait for Clk_period;
		Addr <=  "0100000000100";
		Trees_din <= x"0b008d04";
		wait for Clk_period;
		Addr <=  "0100000000101";
		Trees_din <= x"006820d1";
		wait for Clk_period;
		Addr <=  "0100000000110";
		Trees_din <= x"ffe620d1";
		wait for Clk_period;
		Addr <=  "0100000000111";
		Trees_din <= x"03f67d04";
		wait for Clk_period;
		Addr <=  "0100000001000";
		Trees_din <= x"003720d1";
		wait for Clk_period;
		Addr <=  "0100000001001";
		Trees_din <= x"ff9320d1";
		wait for Clk_period;
		Addr <=  "0100000001010";
		Trees_din <= x"15004c10";
		wait for Clk_period;
		Addr <=  "0100000001011";
		Trees_din <= x"13039808";
		wait for Clk_period;
		Addr <=  "0100000001100";
		Trees_din <= x"13039104";
		wait for Clk_period;
		Addr <=  "0100000001101";
		Trees_din <= x"fffc20d1";
		wait for Clk_period;
		Addr <=  "0100000001110";
		Trees_din <= x"008a20d1";
		wait for Clk_period;
		Addr <=  "0100000001111";
		Trees_din <= x"16006b04";
		wait for Clk_period;
		Addr <=  "0100000010000";
		Trees_din <= x"ff6e20d1";
		wait for Clk_period;
		Addr <=  "0100000010001";
		Trees_din <= x"002c20d1";
		wait for Clk_period;
		Addr <=  "0100000010010";
		Trees_din <= x"10005304";
		wait for Clk_period;
		Addr <=  "0100000010011";
		Trees_din <= x"ff3e20d1";
		wait for Clk_period;
		Addr <=  "0100000010100";
		Trees_din <= x"13027e04";
		wait for Clk_period;
		Addr <=  "0100000010101";
		Trees_din <= x"004e20d1";
		wait for Clk_period;
		Addr <=  "0100000010110";
		Trees_din <= x"ff9a20d1";
		wait for Clk_period;
		Addr <=  "0100000010111";
		Trees_din <= x"1e02762c";
		wait for Clk_period;
		Addr <=  "0100000011000";
		Trees_din <= x"0600931c";
		wait for Clk_period;
		Addr <=  "0100000011001";
		Trees_din <= x"08003b0c";
		wait for Clk_period;
		Addr <=  "0100000011010";
		Trees_din <= x"06ffed08";
		wait for Clk_period;
		Addr <=  "0100000011011";
		Trees_din <= x"05f78604";
		wait for Clk_period;
		Addr <=  "0100000011100";
		Trees_din <= x"008320d1";
		wait for Clk_period;
		Addr <=  "0100000011101";
		Trees_din <= x"ffc820d1";
		wait for Clk_period;
		Addr <=  "0100000011110";
		Trees_din <= x"ff9b20d1";
		wait for Clk_period;
		Addr <=  "0100000011111";
		Trees_din <= x"010ddb08";
		wait for Clk_period;
		Addr <=  "0100000100000";
		Trees_din <= x"04fb2604";
		wait for Clk_period;
		Addr <=  "0100000100001";
		Trees_din <= x"002a20d1";
		wait for Clk_period;
		Addr <=  "0100000100010";
		Trees_din <= x"ff6520d1";
		wait for Clk_period;
		Addr <=  "0100000100011";
		Trees_din <= x"17f71604";
		wait for Clk_period;
		Addr <=  "0100000100100";
		Trees_din <= x"ffc620d1";
		wait for Clk_period;
		Addr <=  "0100000100101";
		Trees_din <= x"007020d1";
		wait for Clk_period;
		Addr <=  "0100000100110";
		Trees_din <= x"08003304";
		wait for Clk_period;
		Addr <=  "0100000100111";
		Trees_din <= x"ffb520d1";
		wait for Clk_period;
		Addr <=  "0100000101000";
		Trees_din <= x"0c007a08";
		wait for Clk_period;
		Addr <=  "0100000101001";
		Trees_din <= x"11003304";
		wait for Clk_period;
		Addr <=  "0100000101010";
		Trees_din <= x"00b220d1";
		wait for Clk_period;
		Addr <=  "0100000101011";
		Trees_din <= x"004220d1";
		wait for Clk_period;
		Addr <=  "0100000101100";
		Trees_din <= x"ffec20d1";
		wait for Clk_period;
		Addr <=  "0100000101101";
		Trees_din <= x"0d02ac0c";
		wait for Clk_period;
		Addr <=  "0100000101110";
		Trees_din <= x"08004404";
		wait for Clk_period;
		Addr <=  "0100000101111";
		Trees_din <= x"00a520d1";
		wait for Clk_period;
		Addr <=  "0100000110000";
		Trees_din <= x"11025904";
		wait for Clk_period;
		Addr <=  "0100000110001";
		Trees_din <= x"005c20d1";
		wait for Clk_period;
		Addr <=  "0100000110010";
		Trees_din <= x"ffe820d1";
		wait for Clk_period;
		Addr <=  "0100000110011";
		Trees_din <= x"ffc720d1";
		wait for Clk_period;
		Addr <=  "0100000110100";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  1
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"000dd180";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"0007a040";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"00055e20";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"05f8ea10";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"02fed208";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"10004604";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"003701a5";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"ff7e01a5";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"17f70004";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"ff9001a5";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"ff5801a5";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"05f90208";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"02050b04";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"ff8c01a5";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"00ca01a5";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"15004204";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"ff6201a5";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"ff9c01a5";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"010ce310";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"02079008";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"08004904";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"fffa01a5";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"017001a5";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"04fd9f04";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"003101a5";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"ff5701a5";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"11000708";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"05f64604";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"ff7401a5";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"015c01a5";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"0b005c04";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"ffae01a5";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"ff5301a5";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"010d1620";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"000b8f10";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"0205d508";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"010a6404";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"027201a5";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"00f001a5";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"04017704";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"00e101a5";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"fffb01a5";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"020b6e08";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"010ab104";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"036a01a5";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"01bf01a5";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"0a003e04";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"015c01a5";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"ffb701a5";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"01100910";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"000c4208";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"07005a04";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"ffc201a5";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"00ca01a5";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"0f000504";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"ffea01a5";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"019601a5";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"0f000008";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"11004904";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"ff9901a5";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"010101a5";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"0d000004";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"002f01a5";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"ff6401a5";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"01102d30";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"000f361c";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"07f6b40c";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"010b2808";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"04051904";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"01f801a5";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"ff9601a5";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"ff7701a5";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"03f4a508";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"010a5104";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"026e01a5";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"ff8c01a5";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"01fed304";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"010201a5";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"038401a5";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"00126b10";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"07f4c808";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"05f36604";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"003701a5";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"015c01a5";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"12009904";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"03f301a5";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"00df01a5";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"04ac01a5";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"01138818";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"00100a0c";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"03f6a108";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"02041804";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"01b701a5";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"002201a5";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"ff6601a5";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"16005b04";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"fff301a5";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"0a004e04";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"02f401a5";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"003701a5";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"1801b908";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"03f5fd04";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"ff5f01a5";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"000001a5";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"005b01a5";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"000b7d78";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"0007a038";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"00055e1c";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"05f8ea0c";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"06fc5f08";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"00036a04";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"ff5e0361";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"ffd90361";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"ff570361";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"0c008508";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"11013704";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"ff820361";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"00f20361";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"00ff8504";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"ff590361";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"ff960361";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"05f5ca10";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"0107ec08";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"1101f804";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"ff740361";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"00d40361";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"0b005c04";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"ffae0361";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"ff590361";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"03fdcb08";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"07fd3804";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"ff8a0361";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"00020361";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"01310361";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"010dac20";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"020a0010";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"010a9f08";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"1101e004";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"015b0361";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"00420361";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"0207cf04";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"009f0361";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"ffc60361";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"05f87508";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"06005504";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"00390361";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"ff5f0361";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"06034b04";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"ff890361";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"014b0361";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"05f55110";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"02027608";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"0c00ab04";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"ff6e0361";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"00610361";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"12007104";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"ffa70361";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"ff5d0361";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"16007308";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"12008c04";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"ff8c0361";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"00a80361";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"08004104";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"018e0361";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"fff50361";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"01107c40";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"000d1b20";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"010d9f10";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"07fbe808";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"02070c04";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"013b0361";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"00730361";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"0403b204";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"01d80361";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"ff7a0361";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"19000008";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"0b005e04";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"011d0361";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"ffa50361";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"11010204";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"01e70361";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"00410361";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"010ea610";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"0c013608";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"0e005304";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"01a10361";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"00bf0361";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"07fb1904";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"00c00361";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"00080361";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"05f4d508";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"06ff5104";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"01860361";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"00c50361";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"08003504";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"00ed0361";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"ff660361";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"00126b1c";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"0f00000c";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"11000a04";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"ff7d0361";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"01147f04";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"01e80361";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"ffa50361";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"000d4108";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"17018904";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"ff6a0361";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"003e0361";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"16005b04";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"ff690361";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"00110361";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"01134408";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"15003704";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"008f0361";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"01d90361";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"ffeb0361";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"000b576c";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"0007a030";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"0003b414";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"13006204";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"002904e5";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"05f99f08";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"02fed204";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"ffc604e5";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"ff5e04e5";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"05f9b704";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"006b04e5";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"ff7e04e5";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"0301e210";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"05f5ca08";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"0107ec04";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"ffce04e5";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"ff6104e5";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"1c026904";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"fffc04e5";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"ff9004e5";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"0e002908";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"1403fb04";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"003304e5";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"020304e5";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"ff8704e5";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"010dac1c";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"04017710";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"05f46508";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"12007304";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"009604e5";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"ff9d04e5";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"16009a04";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"00c904e5";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"ff7104e5";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"16004604";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"018104e5";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"0107b304";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"002e04e5";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"ff8404e5";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"05f55110";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"02076e08";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"02027604";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"ffcd04e5";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"ff6704e5";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"12006f04";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"011d04e5";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"ff6c04e5";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"10004608";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"0b009304";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"ff8504e5";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"007d04e5";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"04fed704";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"011104e5";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"ffb704e5";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"01107c2c";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"0010681c";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"07f5b90c";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"0208e008";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"0206d504";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"ff5c04e5";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"00c504e5";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"ff5404e5";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"010ea608";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"0405f104";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"010304e5";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"002f04e5";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"03f76604";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"00b804e5";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"ffc204e5";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"06f91e04";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"001c04e5";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"1401a208";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"010c7304";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"010304e5";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"fff004e5";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"013504e5";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"00126b1c";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"0f00000c";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"11000a04";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"ff8304e5";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"0111ea04";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"01de04e5";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"003f04e5";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"000d4108";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"17018904";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"ff7004e5";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"00bd04e5";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"0114da04";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"001d04e5";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"ff6c04e5";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"0113440c";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"0e002704";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"001504e5";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"10005104";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"016b04e5";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"007004e5";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"ffee04e5";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"0009cb78";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"0007093c";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"0003b41c";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"05f99f10";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"02fed208";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"03f8cb04";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"004406a9";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"ff9306a9";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"0b005d04";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"ffa906a9";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"ff5e06a9";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"05f9b704";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"006506a9";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"0c008504";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"000a06a9";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"ff7c06a9";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"05f68610";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"0301e208";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"11021c04";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"ff5e06a9";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"ffbd06a9";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"0e002904";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"018806a9";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"ffaa06a9";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"1f026808";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"03f7ad04";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"ff8706a9";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"005006a9";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"21006804";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"ff7d06a9";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"009e06a9";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"010d5f20";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"07fc7110";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"0d010608";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"0b008704";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"ff8206a9";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"006306a9";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"11027a04";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"00b406a9";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"ff7f06a9";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"16006208";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"06ff9c04";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"016306a9";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"004506a9";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"0c009e04";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"00a206a9";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"000006a9";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"1200710c";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"15003c04";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"011a06a9";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"01102d04";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"002c06a9";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"ff6f06a9";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"05f61308";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"06fb1404";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"ffd806a9";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"ff5f06a9";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"0900a604";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"00a106a9";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"ff8506a9";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"01107c34";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"000e8020";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"010e8410";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"07f83c08";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"0a004804";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"007606a9";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"ffaf06a9";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"020bce04";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"00b006a9";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"ffbf06a9";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"06fbd208";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"04ff8604";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"019a06a9";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"002c06a9";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"000c7a04";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"ffa406a9";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"005306a9";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"0e000d04";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"ff8d06a9";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"00126b08";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"04067d04";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"00d806a9";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"003506a9";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"1bfa9c04";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"006a06a9";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"00fc06a9";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"000e1920";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"0f000010";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"0111ea08";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"0b007204";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"001a06a9";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"018f06a9";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"06ffa804";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"ff8b06a9";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"004006a9";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"01112508";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"0d000f04";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"01ab06a9";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"ff9606a9";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"0b006404";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"ffae06a9";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"ff6106a9";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"0114da10";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"0e002608";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"02066904";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"ff7506a9";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"003906a9";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"07f87a04";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"00eb06a9";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"000306a9";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"0c00c804";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"ff7206a9";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"003c06a9";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"0007e660";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"00055e2c";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"02063d20";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"02056b10";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"010ab108";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"0106ed04";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"ff81080d";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"0003080d";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"13011f04";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"0008080d";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"ff6d080d";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"11018108";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"00049604";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"ff71080d";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"002f080d";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"13028c04";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"ff8d080d";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"0124080d";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"17f70a08";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"05f99f04";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"ff7e080d";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"009f080d";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"ff5f080d";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"010c241c";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"02079010";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"0d000b08";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"06fd3704";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"002f080d";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"ff62080d";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"01036904";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"ffa0080d";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"00bd080d";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"04fd9f08";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"1afd4e04";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"00c5080d";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"ff93080d";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"ff5e080d";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"0e003b08";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"05f87504";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"ff61080d";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"0002080d";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"0a004408";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"0f000204";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"0137080d";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"ff9b080d";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"05f2a304";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"0037080d";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"ff70080d";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"000d1b2c";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"010d9f1c";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"04037d10";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"020ad308";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"0c00ac04";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"0055080d";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"009c080d";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"0402ab04";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"ff9c080d";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"00ae080d";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"15003004";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"00ed080d";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"07f80704";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"0046080d";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"ff81080d";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"05f2a304";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"ff63080d";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"08005008";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"18000804";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"0070080d";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"ffd7080d";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"0141080d";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"0113881c";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"00126b10";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"07f65308";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"0d000904";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"ff8c080d";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"0071080d";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"0b007104";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"00c5080d";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"007f080d";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"15001c04";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"0014080d";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"1bfa9c04";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"0059080d";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"00da080d";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"1801b908";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"0900e704";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"ff6e080d";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"0025080d";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"0074080d";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"0007e650";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"0003b428";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"05f99f14";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"02fed208";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"12007604";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"ffa80959";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"00460959";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"0b005d08";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"0c008404";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"ff8a0959";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"00460959";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"ff620959";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"00fe3804";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"ff680959";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"0e003208";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"08004204";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"ff780959";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"001e0959";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"1100dd04";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"ffa50959";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"00760959";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"07fd0414";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"0b005d08";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"0f000604";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"ff8c0959";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"00cc0959";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"14040004";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"ff5f0959";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"15003d04";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"00db0959";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"ff940959";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"01102d10";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"0101e508";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"0007a004";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"ff6b0959";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"00130959";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"0900e204";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"fff10959";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"00680959";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"ff6a0959";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"000fee3c";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"0110b320";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"16009a10";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"000c6908";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"05f37304";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"ffc60959";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"004e0959";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"0405f104";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"007e0959";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"ffbe0959";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"08004608";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"07fa6c04";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"fff40959";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"ff460959";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"17f84804";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"00a70959";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"fff00959";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"0f00000c";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"0c00b008";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"11004704";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"ff7c0959";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"00690959";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"01500959";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"000dd108";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"08004f04";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"ff830959";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"00af0959";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"07f72304";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"ff750959";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"00860959";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"01134414";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"0e000d04";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"ff860959";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"00126b08";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"06fc0304";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"ffe80959";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"009b0959";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"1bfa9c04";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"00470959";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"00c40959";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"0d015304";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"ff7b0959";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"008b0959";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"0007e650";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"00066024";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"02083320";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"010c3410";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"15004108";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"17f70f04";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"006f0abd";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"ff9a0abd";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"0e002d04";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"012e0abd";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"fffc0abd";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"03028708";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"13011f04";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"000d0abd";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"ff640abd";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"04fa6804";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"ff880abd";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"00d00abd";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"ff640abd";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"07fd040c";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"0e003b04";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"ff650abd";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"00c70abd";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"ff870abd";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"0d004810";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"0f000008";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"0a004604";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"010b0abd";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"ff970abd";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"07fdca04";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"00050abd";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"ff740abd";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"1f028408";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"010d5f04";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"00ad0abd";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"ffc30abd";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"17f91b04";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"00140abd";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"ff760abd";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"000fee38";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"0111f820";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"16009a10";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"15004d08";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"01049404";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"008a0abd";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"003a0abd";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"0900d004";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"00fd0abd";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"ff6a0abd";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"08004408";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"08003804";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"ffed0abd";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"ff4b0abd";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"0e005304";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"009e0abd";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"ffca0abd";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"000e190c";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"08003008";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"0c00af04";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"ffac0abd";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"00db0abd";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"ff680abd";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"000e6804";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"010b0abd";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"02042204";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"ff760abd";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"004e0abd";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"00126b1c";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"06fc030c";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"05f34304";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"ff380abd";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"06fb1404";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"00a20abd";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"ffa80abd";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"05f1a608";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"1e028304";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"004b0abd";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"ff440abd";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"04067d04";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"00980abd";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"00020abd";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"0113440c";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"15001c04";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"00010abd";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"0e001b04";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"005f0abd";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"00b40abd";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"00030abd";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"0007e634";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"02088124";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"01102d20";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"00026910";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"0605d608";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"0200d204";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"ffd50bcd";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"ff6e0bcd";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"0a004404";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"00890bcd";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"ff890bcd";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"06feb408";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"05f76d04";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"fff00bcd";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"00b20bcd";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"16007a04";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"ffad0bcd";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"00290bcd";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"ff6a0bcd";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"1400fb04";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"00420bcd";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"1102e204";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"ff640bcd";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"04fd9f04";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"00450bcd";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"ffa40bcd";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"00126b40";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"000c6920";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"05f55d10";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"07fded08";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"10004504";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"00030bcd";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"ffae0bcd";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"03f85204";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"00920bcd";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"ffc50bcd";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"13040008";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"03f91804";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"000e0bcd";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"007a0bcd";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"03f91804";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"014e0bcd";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"fff10bcd";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"04067d10";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"010acf08";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"07f57704";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"ffa10bcd";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"008c0bcd";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"06ff2504";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"005a0bcd";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"00140bcd";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"11015b08";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"00730bcd";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"ff4b0bcd";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"03f61804";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"00a50bcd";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"ffba0bcd";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"15001c04";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"ffff0bcd";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"0113440c";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"0e005308";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"0e001b04";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"004f0bcd";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"00aa0bcd";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"00260bcd";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"00070bcd";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"0007094c";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"02063d2c";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"010b0414";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"00ff8508";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"04fdb904";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"ff6d0d21";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"00000d21";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"0e002404";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"ff750d21";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"15003504";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"01230d21";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"002a0d21";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"0900e208";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"13011f04";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"fffe0d21";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"ff660d21";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"010d7008";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"07000104";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"01610d21";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"ffac0d21";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"14040004";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"ff770d21";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"003c0d21";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"14040010";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"1102d208";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"1e060004";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"ff620d21";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"002f0d21";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"17f80204";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"009d0d21";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"ff850d21";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"10004c0c";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"03f9d108";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"04fdd604";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"018d0d21";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"00200d21";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"ff990d21";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"ff7a0d21";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"00126b38";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"0111f820";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"000b5710";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"05f50308";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"0900ec04";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"ffc70d21";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"007d0d21";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"0f000004";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"00930d21";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"00230d21";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"07f5b908";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"0208ff04";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"00180d21";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"ff3b0d21";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"01066704";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"007f0d21";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"00400d21";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"000e190c";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"08003008";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"0c00af04";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"ffb00d21";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"00bf0d21";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"ff6c0d21";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"12007e08";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"0203b504";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"ffbd0d21";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"00b00d21";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"ff7e0d21";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"010f8d14";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"1f028708";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"01f13b04";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"00050d21";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"00a60d21";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"03f4ba04";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"00920d21";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"0900df04";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"ff470d21";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"005e0d21";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"0900e80c";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"0a004004";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"ffc20d21";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"08004704";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"00b60d21";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"00080d21";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"0204a504";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"ff790d21";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"fffc0d21";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"00070950";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"02063d30";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"010c3418";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"00ff8508";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"04fdb904";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"ff700e55";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"00080e55";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"08004208";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"1403fb04";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"ff8b0e55";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"003f0e55";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"1b026604";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"ff940e55";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"00b20e55";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"03028710";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"00066008";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"13011f04";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"00240e55";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"ff6a0e55";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"05f72704";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"ff8a0e55";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"00ac0e55";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"04fa6804";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"ff9b0e55";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"00c90e55";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"14040010";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"1102d208";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"1e060004";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"ff640e55";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"002d0e55";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"17f80204";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"008a0e55";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"ff8a0e55";
		wait for Clk_period;
		Addr <=  "0001101101001";
		Trees_din <= x"0a00460c";
		wait for Clk_period;
		Addr <=  "0001101101010";
		Trees_din <= x"0c008404";
		wait for Clk_period;
		Addr <=  "0001101101011";
		Trees_din <= x"ff970e55";
		wait for Clk_period;
		Addr <=  "0001101101100";
		Trees_din <= x"17f72c04";
		wait for Clk_period;
		Addr <=  "0001101101101";
		Trees_din <= x"013c0e55";
		wait for Clk_period;
		Addr <=  "0001101101110";
		Trees_din <= x"003b0e55";
		wait for Clk_period;
		Addr <=  "0001101101111";
		Trees_din <= x"ff7f0e55";
		wait for Clk_period;
		Addr <=  "0001101110000";
		Trees_din <= x"00126b24";
		wait for Clk_period;
		Addr <=  "0001101110001";
		Trees_din <= x"0114da20";
		wait for Clk_period;
		Addr <=  "0001101110010";
		Trees_din <= x"000c6910";
		wait for Clk_period;
		Addr <=  "0001101110011";
		Trees_din <= x"07fcbd08";
		wait for Clk_period;
		Addr <=  "0001101110100";
		Trees_din <= x"0a004e04";
		wait for Clk_period;
		Addr <=  "0001101110101";
		Trees_din <= x"ffea0e55";
		wait for Clk_period;
		Addr <=  "0001101110110";
		Trees_din <= x"00620e55";
		wait for Clk_period;
		Addr <=  "0001101110111";
		Trees_din <= x"1e028504";
		wait for Clk_period;
		Addr <=  "0001101111000";
		Trees_din <= x"004d0e55";
		wait for Clk_period;
		Addr <=  "0001101111001";
		Trees_din <= x"ffce0e55";
		wait for Clk_period;
		Addr <=  "0001101111010";
		Trees_din <= x"04067d08";
		wait for Clk_period;
		Addr <=  "0001101111011";
		Trees_din <= x"01066704";
		wait for Clk_period;
		Addr <=  "0001101111100";
		Trees_din <= x"008a0e55";
		wait for Clk_period;
		Addr <=  "0001101111101";
		Trees_din <= x"00360e55";
		wait for Clk_period;
		Addr <=  "0001101111110";
		Trees_din <= x"11015b04";
		wait for Clk_period;
		Addr <=  "0001101111111";
		Trees_din <= x"ff8a0e55";
		wait for Clk_period;
		Addr <=  "0001110000000";
		Trees_din <= x"002d0e55";
		wait for Clk_period;
		Addr <=  "0001110000001";
		Trees_din <= x"ff790e55";
		wait for Clk_period;
		Addr <=  "0001110000010";
		Trees_din <= x"010f8d14";
		wait for Clk_period;
		Addr <=  "0001110000011";
		Trees_din <= x"1f02870c";
		wait for Clk_period;
		Addr <=  "0001110000100";
		Trees_din <= x"01f13b04";
		wait for Clk_period;
		Addr <=  "0001110000101";
		Trees_din <= x"00020e55";
		wait for Clk_period;
		Addr <=  "0001110000110";
		Trees_din <= x"05f0b704";
		wait for Clk_period;
		Addr <=  "0001110000111";
		Trees_din <= x"00550e55";
		wait for Clk_period;
		Addr <=  "0001110001000";
		Trees_din <= x"00a30e55";
		wait for Clk_period;
		Addr <=  "0001110001001";
		Trees_din <= x"03f4ba04";
		wait for Clk_period;
		Addr <=  "0001110001010";
		Trees_din <= x"00870e55";
		wait for Clk_period;
		Addr <=  "0001110001011";
		Trees_din <= x"ffc20e55";
		wait for Clk_period;
		Addr <=  "0001110001100";
		Trees_din <= x"0900e80c";
		wait for Clk_period;
		Addr <=  "0001110001101";
		Trees_din <= x"07f80708";
		wait for Clk_period;
		Addr <=  "0001110001110";
		Trees_din <= x"0e004104";
		wait for Clk_period;
		Addr <=  "0001110001111";
		Trees_din <= x"00af0e55";
		wait for Clk_period;
		Addr <=  "0001110010000";
		Trees_din <= x"00010e55";
		wait for Clk_period;
		Addr <=  "0001110010001";
		Trees_din <= x"ffc80e55";
		wait for Clk_period;
		Addr <=  "0001110010010";
		Trees_din <= x"0b006404";
		wait for Clk_period;
		Addr <=  "0001110010011";
		Trees_din <= x"00630e55";
		wait for Clk_period;
		Addr <=  "0001110010100";
		Trees_din <= x"ff3a0e55";
		wait for Clk_period;
		Addr <=  "0001110010101";
		Trees_din <= x"0009b250";
		wait for Clk_period;
		Addr <=  "0001110010110";
		Trees_din <= x"0003b428";
		wait for Clk_period;
		Addr <=  "0001110010111";
		Trees_din <= x"0200d210";
		wait for Clk_period;
		Addr <=  "0001110011000";
		Trees_din <= x"04f98804";
		wait for Clk_period;
		Addr <=  "0001110011001";
		Trees_din <= x"ff850f71";
		wait for Clk_period;
		Addr <=  "0001110011010";
		Trees_din <= x"1afcf808";
		wait for Clk_period;
		Addr <=  "0001110011011";
		Trees_din <= x"1100e504";
		wait for Clk_period;
		Addr <=  "0001110011100";
		Trees_din <= x"01530f71";
		wait for Clk_period;
		Addr <=  "0001110011101";
		Trees_din <= x"00150f71";
		wait for Clk_period;
		Addr <=  "0001110011110";
		Trees_din <= x"ff970f71";
		wait for Clk_period;
		Addr <=  "0001110011111";
		Trees_din <= x"0e00390c";
		wait for Clk_period;
		Addr <=  "0001110100000";
		Trees_din <= x"16004808";
		wait for Clk_period;
		Addr <=  "0001110100001";
		Trees_din <= x"0d01b204";
		wait for Clk_period;
		Addr <=  "0001110100010";
		Trees_din <= x"ffa40f71";
		wait for Clk_period;
		Addr <=  "0001110100011";
		Trees_din <= x"00400f71";
		wait for Clk_period;
		Addr <=  "0001110100100";
		Trees_din <= x"ff660f71";
		wait for Clk_period;
		Addr <=  "0001110100101";
		Trees_din <= x"0e003a04";
		wait for Clk_period;
		Addr <=  "0001110100110";
		Trees_din <= x"00ea0f71";
		wait for Clk_period;
		Addr <=  "0001110100111";
		Trees_din <= x"19000404";
		wait for Clk_period;
		Addr <=  "0001110101000";
		Trees_din <= x"ff960f71";
		wait for Clk_period;
		Addr <=  "0001110101001";
		Trees_din <= x"00750f71";
		wait for Clk_period;
		Addr <=  "0001110101010";
		Trees_din <= x"05f38308";
		wait for Clk_period;
		Addr <=  "0001110101011";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0001110101100";
		Trees_din <= x"00840f71";
		wait for Clk_period;
		Addr <=  "0001110101101";
		Trees_din <= x"ff640f71";
		wait for Clk_period;
		Addr <=  "0001110101110";
		Trees_din <= x"04fde910";
		wait for Clk_period;
		Addr <=  "0001110101111";
		Trees_din <= x"15003708";
		wait for Clk_period;
		Addr <=  "0001110110000";
		Trees_din <= x"06ff1504";
		wait for Clk_period;
		Addr <=  "0001110110001";
		Trees_din <= x"00c40f71";
		wait for Clk_period;
		Addr <=  "0001110110010";
		Trees_din <= x"00000f71";
		wait for Clk_period;
		Addr <=  "0001110110011";
		Trees_din <= x"0b006004";
		wait for Clk_period;
		Addr <=  "0001110110100";
		Trees_din <= x"009a0f71";
		wait for Clk_period;
		Addr <=  "0001110110101";
		Trees_din <= x"fff10f71";
		wait for Clk_period;
		Addr <=  "0001110110110";
		Trees_din <= x"08003d08";
		wait for Clk_period;
		Addr <=  "0001110110111";
		Trees_din <= x"08003904";
		wait for Clk_period;
		Addr <=  "0001110111000";
		Trees_din <= x"ffd30f71";
		wait for Clk_period;
		Addr <=  "0001110111001";
		Trees_din <= x"ff570f71";
		wait for Clk_period;
		Addr <=  "0001110111010";
		Trees_din <= x"03f87d04";
		wait for Clk_period;
		Addr <=  "0001110111011";
		Trees_din <= x"ffc70f71";
		wait for Clk_period;
		Addr <=  "0001110111100";
		Trees_din <= x"003a0f71";
		wait for Clk_period;
		Addr <=  "0001110111101";
		Trees_din <= x"0012e528";
		wait for Clk_period;
		Addr <=  "0001110111110";
		Trees_din <= x"020eae20";
		wait for Clk_period;
		Addr <=  "0001110111111";
		Trees_din <= x"0105ad10";
		wait for Clk_period;
		Addr <=  "0001111000000";
		Trees_din <= x"1c023a08";
		wait for Clk_period;
		Addr <=  "0001111000001";
		Trees_din <= x"02082604";
		wait for Clk_period;
		Addr <=  "0001111000010";
		Trees_din <= x"ff3c0f71";
		wait for Clk_period;
		Addr <=  "0001111000011";
		Trees_din <= x"00140f71";
		wait for Clk_period;
		Addr <=  "0001111000100";
		Trees_din <= x"0b007b04";
		wait for Clk_period;
		Addr <=  "0001111000101";
		Trees_din <= x"009d0f71";
		wait for Clk_period;
		Addr <=  "0001111000110";
		Trees_din <= x"001e0f71";
		wait for Clk_period;
		Addr <=  "0001111000111";
		Trees_din <= x"020a3108";
		wait for Clk_period;
		Addr <=  "0001111001000";
		Trees_din <= x"16009604";
		wait for Clk_period;
		Addr <=  "0001111001001";
		Trees_din <= x"00300f71";
		wait for Clk_period;
		Addr <=  "0001111001010";
		Trees_din <= x"ffcd0f71";
		wait for Clk_period;
		Addr <=  "0001111001011";
		Trees_din <= x"0b007104";
		wait for Clk_period;
		Addr <=  "0001111001100";
		Trees_din <= x"ff500f71";
		wait for Clk_period;
		Addr <=  "0001111001101";
		Trees_din <= x"000e0f71";
		wait for Clk_period;
		Addr <=  "0001111001110";
		Trees_din <= x"05f4c304";
		wait for Clk_period;
		Addr <=  "0001111001111";
		Trees_din <= x"ffe90f71";
		wait for Clk_period;
		Addr <=  "0001111010000";
		Trees_din <= x"ff590f71";
		wait for Clk_period;
		Addr <=  "0001111010001";
		Trees_din <= x"0e001c0c";
		wait for Clk_period;
		Addr <=  "0001111010010";
		Trees_din <= x"0e001a08";
		wait for Clk_period;
		Addr <=  "0001111010011";
		Trees_din <= x"15001c04";
		wait for Clk_period;
		Addr <=  "0001111010100";
		Trees_din <= x"fff00f71";
		wait for Clk_period;
		Addr <=  "0001111010101";
		Trees_din <= x"007b0f71";
		wait for Clk_period;
		Addr <=  "0001111010110";
		Trees_din <= x"ff810f71";
		wait for Clk_period;
		Addr <=  "0001111010111";
		Trees_din <= x"1803a108";
		wait for Clk_period;
		Addr <=  "0001111011000";
		Trees_din <= x"01134404";
		wait for Clk_period;
		Addr <=  "0001111011001";
		Trees_din <= x"00980f71";
		wait for Clk_period;
		Addr <=  "0001111011010";
		Trees_din <= x"001a0f71";
		wait for Clk_period;
		Addr <=  "0001111011011";
		Trees_din <= x"fffb0f71";
		wait for Clk_period;
		Addr <=  "0001111011100";
		Trees_din <= x"0007092c";
		wait for Clk_period;
		Addr <=  "0001111011101";
		Trees_din <= x"1f028428";
		wait for Clk_period;
		Addr <=  "0001111011110";
		Trees_din <= x"04000320";
		wait for Clk_period;
		Addr <=  "0001111011111";
		Trees_din <= x"05f76110";
		wait for Clk_period;
		Addr <=  "0001111100000";
		Trees_din <= x"11018e08";
		wait for Clk_period;
		Addr <=  "0001111100001";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0001111100010";
		Trees_din <= x"00041035";
		wait for Clk_period;
		Addr <=  "0001111100011";
		Trees_din <= x"ff7a1035";
		wait for Clk_period;
		Addr <=  "0001111100100";
		Trees_din <= x"13032e04";
		wait for Clk_period;
		Addr <=  "0001111100101";
		Trees_din <= x"ffe31035";
		wait for Clk_period;
		Addr <=  "0001111100110";
		Trees_din <= x"00921035";
		wait for Clk_period;
		Addr <=  "0001111100111";
		Trees_din <= x"00055e08";
		wait for Clk_period;
		Addr <=  "0001111101000";
		Trees_din <= x"0b008804";
		wait for Clk_period;
		Addr <=  "0001111101001";
		Trees_din <= x"00061035";
		wait for Clk_period;
		Addr <=  "0001111101010";
		Trees_din <= x"ff781035";
		wait for Clk_period;
		Addr <=  "0001111101011";
		Trees_din <= x"07036e04";
		wait for Clk_period;
		Addr <=  "0001111101100";
		Trees_din <= x"00b51035";
		wait for Clk_period;
		Addr <=  "0001111101101";
		Trees_din <= x"ff9a1035";
		wait for Clk_period;
		Addr <=  "0001111101110";
		Trees_din <= x"1b037604";
		wait for Clk_period;
		Addr <=  "0001111101111";
		Trees_din <= x"ff6a1035";
		wait for Clk_period;
		Addr <=  "0001111110000";
		Trees_din <= x"00201035";
		wait for Clk_period;
		Addr <=  "0001111110001";
		Trees_din <= x"ff6b1035";
		wait for Clk_period;
		Addr <=  "0001111110010";
		Trees_din <= x"0012e520";
		wait for Clk_period;
		Addr <=  "0001111110011";
		Trees_din <= x"01f76408";
		wait for Clk_period;
		Addr <=  "0001111110100";
		Trees_din <= x"0900b304";
		wait for Clk_period;
		Addr <=  "0001111110101";
		Trees_din <= x"003c1035";
		wait for Clk_period;
		Addr <=  "0001111110110";
		Trees_din <= x"ff441035";
		wait for Clk_period;
		Addr <=  "0001111110111";
		Trees_din <= x"1c02880c";
		wait for Clk_period;
		Addr <=  "0001111111000";
		Trees_din <= x"0114da08";
		wait for Clk_period;
		Addr <=  "0001111111001";
		Trees_din <= x"02020604";
		wait for Clk_period;
		Addr <=  "0001111111010";
		Trees_din <= x"00731035";
		wait for Clk_period;
		Addr <=  "0001111111011";
		Trees_din <= x"00211035";
		wait for Clk_period;
		Addr <=  "0001111111100";
		Trees_din <= x"ff811035";
		wait for Clk_period;
		Addr <=  "0001111111101";
		Trees_din <= x"1e028808";
		wait for Clk_period;
		Addr <=  "0001111111110";
		Trees_din <= x"1400fb04";
		wait for Clk_period;
		Addr <=  "0001111111111";
		Trees_din <= x"00121035";
		wait for Clk_period;
		Addr <=  "0010000000000";
		Trees_din <= x"ff5b1035";
		wait for Clk_period;
		Addr <=  "0010000000001";
		Trees_din <= x"005b1035";
		wait for Clk_period;
		Addr <=  "0010000000010";
		Trees_din <= x"0e001c08";
		wait for Clk_period;
		Addr <=  "0010000000011";
		Trees_din <= x"0014ec04";
		wait for Clk_period;
		Addr <=  "0010000000100";
		Trees_din <= x"ffa81035";
		wait for Clk_period;
		Addr <=  "0010000000101";
		Trees_din <= x"00661035";
		wait for Clk_period;
		Addr <=  "0010000000110";
		Trees_din <= x"1803a10c";
		wait for Clk_period;
		Addr <=  "0010000000111";
		Trees_din <= x"010c8404";
		wait for Clk_period;
		Addr <=  "0010000001000";
		Trees_din <= x"009f1035";
		wait for Clk_period;
		Addr <=  "0010000001001";
		Trees_din <= x"06004f04";
		wait for Clk_period;
		Addr <=  "0010000001010";
		Trees_din <= x"00861035";
		wait for Clk_period;
		Addr <=  "0010000001011";
		Trees_din <= x"ffbf1035";
		wait for Clk_period;
		Addr <=  "0010000001100";
		Trees_din <= x"fffa1035";
		wait for Clk_period;
		Addr <=  "0010000001101";
		Trees_din <= x"00062634";
		wait for Clk_period;
		Addr <=  "0010000001110";
		Trees_din <= x"02083330";
		wait for Clk_period;
		Addr <=  "0010000001111";
		Trees_din <= x"17f71614";
		wait for Clk_period;
		Addr <=  "0010000010000";
		Trees_din <= x"04fc3708";
		wait for Clk_period;
		Addr <=  "0010000010001";
		Trees_din <= x"03033e04";
		wait for Clk_period;
		Addr <=  "0010000010010";
		Trees_din <= x"ff8e1149";
		wait for Clk_period;
		Addr <=  "0010000010011";
		Trees_din <= x"00151149";
		wait for Clk_period;
		Addr <=  "0010000010100";
		Trees_din <= x"0a004608";
		wait for Clk_period;
		Addr <=  "0010000010101";
		Trees_din <= x"0b006d04";
		wait for Clk_period;
		Addr <=  "0010000010110";
		Trees_din <= x"005a1149";
		wait for Clk_period;
		Addr <=  "0010000010111";
		Trees_din <= x"01381149";
		wait for Clk_period;
		Addr <=  "0010000011000";
		Trees_din <= x"fffe1149";
		wait for Clk_period;
		Addr <=  "0010000011001";
		Trees_din <= x"05f8660c";
		wait for Clk_period;
		Addr <=  "0010000011010";
		Trees_din <= x"06fc5f08";
		wait for Clk_period;
		Addr <=  "0010000011011";
		Trees_din <= x"07002004";
		wait for Clk_period;
		Addr <=  "0010000011100";
		Trees_din <= x"00b41149";
		wait for Clk_period;
		Addr <=  "0010000011101";
		Trees_din <= x"ffc31149";
		wait for Clk_period;
		Addr <=  "0010000011110";
		Trees_din <= x"ff671149";
		wait for Clk_period;
		Addr <=  "0010000011111";
		Trees_din <= x"15004108";
		wait for Clk_period;
		Addr <=  "0010000100000";
		Trees_din <= x"0c00ba04";
		wait for Clk_period;
		Addr <=  "0010000100001";
		Trees_din <= x"ff951149";
		wait for Clk_period;
		Addr <=  "0010000100010";
		Trees_din <= x"00191149";
		wait for Clk_period;
		Addr <=  "0010000100011";
		Trees_din <= x"15004704";
		wait for Clk_period;
		Addr <=  "0010000100100";
		Trees_din <= x"009f1149";
		wait for Clk_period;
		Addr <=  "0010000100101";
		Trees_din <= x"ffca1149";
		wait for Clk_period;
		Addr <=  "0010000100110";
		Trees_din <= x"ff6f1149";
		wait for Clk_period;
		Addr <=  "0010000100111";
		Trees_din <= x"0012e53c";
		wait for Clk_period;
		Addr <=  "0010000101000";
		Trees_din <= x"12005d1c";
		wait for Clk_period;
		Addr <=  "0010000101001";
		Trees_din <= x"0a003f0c";
		wait for Clk_period;
		Addr <=  "0010000101010";
		Trees_din <= x"11000404";
		wait for Clk_period;
		Addr <=  "0010000101011";
		Trees_din <= x"ffa11149";
		wait for Clk_period;
		Addr <=  "0010000101100";
		Trees_din <= x"0f000104";
		wait for Clk_period;
		Addr <=  "0010000101101";
		Trees_din <= x"00c21149";
		wait for Clk_period;
		Addr <=  "0010000101110";
		Trees_din <= x"ffb71149";
		wait for Clk_period;
		Addr <=  "0010000101111";
		Trees_din <= x"06ff1a08";
		wait for Clk_period;
		Addr <=  "0010000110000";
		Trees_din <= x"0900cf04";
		wait for Clk_period;
		Addr <=  "0010000110001";
		Trees_din <= x"ff6e1149";
		wait for Clk_period;
		Addr <=  "0010000110010";
		Trees_din <= x"00301149";
		wait for Clk_period;
		Addr <=  "0010000110011";
		Trees_din <= x"04032304";
		wait for Clk_period;
		Addr <=  "0010000110100";
		Trees_din <= x"ff451149";
		wait for Clk_period;
		Addr <=  "0010000110101";
		Trees_din <= x"ffc31149";
		wait for Clk_period;
		Addr <=  "0010000110110";
		Trees_din <= x"13040010";
		wait for Clk_period;
		Addr <=  "0010000110111";
		Trees_din <= x"0e003f08";
		wait for Clk_period;
		Addr <=  "0010000111000";
		Trees_din <= x"10004d04";
		wait for Clk_period;
		Addr <=  "0010000111001";
		Trees_din <= x"00181149";
		wait for Clk_period;
		Addr <=  "0010000111010";
		Trees_din <= x"ffde1149";
		wait for Clk_period;
		Addr <=  "0010000111011";
		Trees_din <= x"000aa704";
		wait for Clk_period;
		Addr <=  "0010000111100";
		Trees_din <= x"fffd1149";
		wait for Clk_period;
		Addr <=  "0010000111101";
		Trees_din <= x"006c1149";
		wait for Clk_period;
		Addr <=  "0010000111110";
		Trees_din <= x"06008908";
		wait for Clk_period;
		Addr <=  "0010000111111";
		Trees_din <= x"12007a04";
		wait for Clk_period;
		Addr <=  "0010001000000";
		Trees_din <= x"01141149";
		wait for Clk_period;
		Addr <=  "0010001000001";
		Trees_din <= x"00351149";
		wait for Clk_period;
		Addr <=  "0010001000010";
		Trees_din <= x"1afd4904";
		wait for Clk_period;
		Addr <=  "0010001000011";
		Trees_din <= x"ff8f1149";
		wait for Clk_period;
		Addr <=  "0010001000100";
		Trees_din <= x"00591149";
		wait for Clk_period;
		Addr <=  "0010001000101";
		Trees_din <= x"0e001c0c";
		wait for Clk_period;
		Addr <=  "0010001000110";
		Trees_din <= x"0e001a08";
		wait for Clk_period;
		Addr <=  "0010001000111";
		Trees_din <= x"0a003204";
		wait for Clk_period;
		Addr <=  "0010001001000";
		Trees_din <= x"ffec1149";
		wait for Clk_period;
		Addr <=  "0010001001001";
		Trees_din <= x"006e1149";
		wait for Clk_period;
		Addr <=  "0010001001010";
		Trees_din <= x"ff8f1149";
		wait for Clk_period;
		Addr <=  "0010001001011";
		Trees_din <= x"1803a10c";
		wait for Clk_period;
		Addr <=  "0010001001100";
		Trees_din <= x"010c8404";
		wait for Clk_period;
		Addr <=  "0010001001101";
		Trees_din <= x"009c1149";
		wait for Clk_period;
		Addr <=  "0010001001110";
		Trees_din <= x"06004f04";
		wait for Clk_period;
		Addr <=  "0010001001111";
		Trees_din <= x"007e1149";
		wait for Clk_period;
		Addr <=  "0010001010000";
		Trees_din <= x"ffc11149";
		wait for Clk_period;
		Addr <=  "0010001010001";
		Trees_din <= x"fff31149";
		wait for Clk_period;
		Addr <=  "0010001010010";
		Trees_din <= x"00126b64";
		wait for Clk_period;
		Addr <=  "0010001010011";
		Trees_din <= x"00062624";
		wait for Clk_period;
		Addr <=  "0010001010100";
		Trees_din <= x"04fdfc14";
		wait for Clk_period;
		Addr <=  "0010001010101";
		Trees_din <= x"17f8f510";
		wait for Clk_period;
		Addr <=  "0010001010110";
		Trees_din <= x"05fb6b08";
		wait for Clk_period;
		Addr <=  "0010001010111";
		Trees_din <= x"1403f504";
		wait for Clk_period;
		Addr <=  "0010001011000";
		Trees_din <= x"ff891255";
		wait for Clk_period;
		Addr <=  "0010001011001";
		Trees_din <= x"00051255";
		wait for Clk_period;
		Addr <=  "0010001011010";
		Trees_din <= x"05ffdc04";
		wait for Clk_period;
		Addr <=  "0010001011011";
		Trees_din <= x"00ab1255";
		wait for Clk_period;
		Addr <=  "0010001011100";
		Trees_din <= x"ffea1255";
		wait for Clk_period;
		Addr <=  "0010001011101";
		Trees_din <= x"ff721255";
		wait for Clk_period;
		Addr <=  "0010001011110";
		Trees_din <= x"1c023c08";
		wait for Clk_period;
		Addr <=  "0010001011111";
		Trees_din <= x"10004904";
		wait for Clk_period;
		Addr <=  "0010001100000";
		Trees_din <= x"00081255";
		wait for Clk_period;
		Addr <=  "0010001100001";
		Trees_din <= x"00251255";
		wait for Clk_period;
		Addr <=  "0010001100010";
		Trees_din <= x"0a005904";
		wait for Clk_period;
		Addr <=  "0010001100011";
		Trees_din <= x"ff6a1255";
		wait for Clk_period;
		Addr <=  "0010001100100";
		Trees_din <= x"000a1255";
		wait for Clk_period;
		Addr <=  "0010001100101";
		Trees_din <= x"04020720";
		wait for Clk_period;
		Addr <=  "0010001100110";
		Trees_din <= x"020ad310";
		wait for Clk_period;
		Addr <=  "0010001100111";
		Trees_din <= x"1b073c08";
		wait for Clk_period;
		Addr <=  "0010001101000";
		Trees_din <= x"0f00f104";
		wait for Clk_period;
		Addr <=  "0010001101001";
		Trees_din <= x"00271255";
		wait for Clk_period;
		Addr <=  "0010001101010";
		Trees_din <= x"ffe91255";
		wait for Clk_period;
		Addr <=  "0010001101011";
		Trees_din <= x"0a004804";
		wait for Clk_period;
		Addr <=  "0010001101100";
		Trees_din <= x"00f31255";
		wait for Clk_period;
		Addr <=  "0010001101101";
		Trees_din <= x"00221255";
		wait for Clk_period;
		Addr <=  "0010001101110";
		Trees_din <= x"12008408";
		wait for Clk_period;
		Addr <=  "0010001101111";
		Trees_din <= x"000d8e04";
		wait for Clk_period;
		Addr <=  "0010001110000";
		Trees_din <= x"ff641255";
		wait for Clk_period;
		Addr <=  "0010001110001";
		Trees_din <= x"fff71255";
		wait for Clk_period;
		Addr <=  "0010001110010";
		Trees_din <= x"01036904";
		wait for Clk_period;
		Addr <=  "0010001110011";
		Trees_din <= x"00991255";
		wait for Clk_period;
		Addr <=  "0010001110100";
		Trees_din <= x"ffdf1255";
		wait for Clk_period;
		Addr <=  "0010001110101";
		Trees_din <= x"0601f910";
		wait for Clk_period;
		Addr <=  "0010001110110";
		Trees_din <= x"1afa7508";
		wait for Clk_period;
		Addr <=  "0010001110111";
		Trees_din <= x"1102d804";
		wait for Clk_period;
		Addr <=  "0010001111000";
		Trees_din <= x"00911255";
		wait for Clk_period;
		Addr <=  "0010001111001";
		Trees_din <= x"ffc21255";
		wait for Clk_period;
		Addr <=  "0010001111010";
		Trees_din <= x"0a004304";
		wait for Clk_period;
		Addr <=  "0010001111011";
		Trees_din <= x"ffa31255";
		wait for Clk_period;
		Addr <=  "0010001111100";
		Trees_din <= x"00011255";
		wait for Clk_period;
		Addr <=  "0010001111101";
		Trees_din <= x"17f7a108";
		wait for Clk_period;
		Addr <=  "0010001111110";
		Trees_din <= x"1e024f04";
		wait for Clk_period;
		Addr <=  "0010001111111";
		Trees_din <= x"fff01255";
		wait for Clk_period;
		Addr <=  "0010010000000";
		Trees_din <= x"00ce1255";
		wait for Clk_period;
		Addr <=  "0010010000001";
		Trees_din <= x"0a004104";
		wait for Clk_period;
		Addr <=  "0010010000010";
		Trees_din <= x"006e1255";
		wait for Clk_period;
		Addr <=  "0010010000011";
		Trees_din <= x"ff931255";
		wait for Clk_period;
		Addr <=  "0010010000100";
		Trees_din <= x"0016b420";
		wait for Clk_period;
		Addr <=  "0010010000101";
		Trees_din <= x"02089614";
		wait for Clk_period;
		Addr <=  "0010010000110";
		Trees_din <= x"010f8d08";
		wait for Clk_period;
		Addr <=  "0010010000111";
		Trees_din <= x"06fb8b04";
		wait for Clk_period;
		Addr <=  "0010010001000";
		Trees_din <= x"000c1255";
		wait for Clk_period;
		Addr <=  "0010010001001";
		Trees_din <= x"00971255";
		wait for Clk_period;
		Addr <=  "0010010001010";
		Trees_din <= x"0900e808";
		wait for Clk_period;
		Addr <=  "0010010001011";
		Trees_din <= x"0b006804";
		wait for Clk_period;
		Addr <=  "0010010001100";
		Trees_din <= x"ffde1255";
		wait for Clk_period;
		Addr <=  "0010010001101";
		Trees_din <= x"006f1255";
		wait for Clk_period;
		Addr <=  "0010010001110";
		Trees_din <= x"ff6f1255";
		wait for Clk_period;
		Addr <=  "0010010001111";
		Trees_din <= x"0108e508";
		wait for Clk_period;
		Addr <=  "0010010010000";
		Trees_din <= x"08003304";
		wait for Clk_period;
		Addr <=  "0010010010001";
		Trees_din <= x"ffe71255";
		wait for Clk_period;
		Addr <=  "0010010010010";
		Trees_din <= x"007c1255";
		wait for Clk_period;
		Addr <=  "0010010010011";
		Trees_din <= x"ff2e1255";
		wait for Clk_period;
		Addr <=  "0010010010100";
		Trees_din <= x"009a1255";
		wait for Clk_period;
		Addr <=  "0010010010101";
		Trees_din <= x"0012e548";
		wait for Clk_period;
		Addr <=  "0010010010110";
		Trees_din <= x"0003b424";
		wait for Clk_period;
		Addr <=  "0010010010111";
		Trees_din <= x"0200d210";
		wait for Clk_period;
		Addr <=  "0010010011000";
		Trees_din <= x"10004b0c";
		wait for Clk_period;
		Addr <=  "0010010011001";
		Trees_din <= x"04f98804";
		wait for Clk_period;
		Addr <=  "0010010011010";
		Trees_din <= x"ffa51321";
		wait for Clk_period;
		Addr <=  "0010010011011";
		Trees_din <= x"1afc5404";
		wait for Clk_period;
		Addr <=  "0010010011100";
		Trees_din <= x"00f51321";
		wait for Clk_period;
		Addr <=  "0010010011101";
		Trees_din <= x"00001321";
		wait for Clk_period;
		Addr <=  "0010010011110";
		Trees_din <= x"ff8e1321";
		wait for Clk_period;
		Addr <=  "0010010011111";
		Trees_din <= x"0e003908";
		wait for Clk_period;
		Addr <=  "0010010100000";
		Trees_din <= x"03f5e504";
		wait for Clk_period;
		Addr <=  "0010010100001";
		Trees_din <= x"00021321";
		wait for Clk_period;
		Addr <=  "0010010100010";
		Trees_din <= x"ff6a1321";
		wait for Clk_period;
		Addr <=  "0010010100011";
		Trees_din <= x"0e003a04";
		wait for Clk_period;
		Addr <=  "0010010100100";
		Trees_din <= x"00ad1321";
		wait for Clk_period;
		Addr <=  "0010010100101";
		Trees_din <= x"07fff404";
		wait for Clk_period;
		Addr <=  "0010010100110";
		Trees_din <= x"002a1321";
		wait for Clk_period;
		Addr <=  "0010010100111";
		Trees_din <= x"ff7e1321";
		wait for Clk_period;
		Addr <=  "0010010101000";
		Trees_din <= x"07097920";
		wait for Clk_period;
		Addr <=  "0010010101001";
		Trees_din <= x"00041110";
		wait for Clk_period;
		Addr <=  "0010010101010";
		Trees_din <= x"06feb408";
		wait for Clk_period;
		Addr <=  "0010010101011";
		Trees_din <= x"0a004404";
		wait for Clk_period;
		Addr <=  "0010010101100";
		Trees_din <= x"019a1321";
		wait for Clk_period;
		Addr <=  "0010010101101";
		Trees_din <= x"001b1321";
		wait for Clk_period;
		Addr <=  "0010010101110";
		Trees_din <= x"1c026204";
		wait for Clk_period;
		Addr <=  "0010010101111";
		Trees_din <= x"00201321";
		wait for Clk_period;
		Addr <=  "0010010110000";
		Trees_din <= x"ffa81321";
		wait for Clk_period;
		Addr <=  "0010010110001";
		Trees_din <= x"0009b208";
		wait for Clk_period;
		Addr <=  "0010010110010";
		Trees_din <= x"07f8a004";
		wait for Clk_period;
		Addr <=  "0010010110011";
		Trees_din <= x"ff801321";
		wait for Clk_period;
		Addr <=  "0010010110100";
		Trees_din <= x"00021321";
		wait for Clk_period;
		Addr <=  "0010010110101";
		Trees_din <= x"06fc5f04";
		wait for Clk_period;
		Addr <=  "0010010110110";
		Trees_din <= x"ffda1321";
		wait for Clk_period;
		Addr <=  "0010010110111";
		Trees_din <= x"001e1321";
		wait for Clk_period;
		Addr <=  "0010010111000";
		Trees_din <= x"ff5e1321";
		wait for Clk_period;
		Addr <=  "0010010111001";
		Trees_din <= x"0e001c08";
		wait for Clk_period;
		Addr <=  "0010010111010";
		Trees_din <= x"0014ec04";
		wait for Clk_period;
		Addr <=  "0010010111011";
		Trees_din <= x"ffa91321";
		wait for Clk_period;
		Addr <=  "0010010111100";
		Trees_din <= x"004b1321";
		wait for Clk_period;
		Addr <=  "0010010111101";
		Trees_din <= x"1803a114";
		wait for Clk_period;
		Addr <=  "0010010111110";
		Trees_din <= x"010c8404";
		wait for Clk_period;
		Addr <=  "0010010111111";
		Trees_din <= x"00961321";
		wait for Clk_period;
		Addr <=  "0010011000000";
		Trees_din <= x"06004f08";
		wait for Clk_period;
		Addr <=  "0010011000001";
		Trees_din <= x"0111c204";
		wait for Clk_period;
		Addr <=  "0010011000010";
		Trees_din <= x"008e1321";
		wait for Clk_period;
		Addr <=  "0010011000011";
		Trees_din <= x"00231321";
		wait for Clk_period;
		Addr <=  "0010011000100";
		Trees_din <= x"00153704";
		wait for Clk_period;
		Addr <=  "0010011000101";
		Trees_din <= x"00551321";
		wait for Clk_period;
		Addr <=  "0010011000110";
		Trees_din <= x"ff601321";
		wait for Clk_period;
		Addr <=  "0010011000111";
		Trees_din <= x"ffe81321";
		wait for Clk_period;
		Addr <=  "0010011001000";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0010011001001";
		Trees_din <= x"0016b474";
		wait for Clk_period;
		Addr <=  "0010011001010";
		Trees_din <= x"0007e638";
		wait for Clk_period;
		Addr <=  "0010011001011";
		Trees_din <= x"0b007e1c";
		wait for Clk_period;
		Addr <=  "0010011001100";
		Trees_din <= x"0b007b0c";
		wait for Clk_period;
		Addr <=  "0010011001101";
		Trees_din <= x"1c028408";
		wait for Clk_period;
		Addr <=  "0010011001110";
		Trees_din <= x"13039604";
		wait for Clk_period;
		Addr <=  "0010011001111";
		Trees_din <= x"00361419";
		wait for Clk_period;
		Addr <=  "0010011010000";
		Trees_din <= x"ffd71419";
		wait for Clk_period;
		Addr <=  "0010011010001";
		Trees_din <= x"ff721419";
		wait for Clk_period;
		Addr <=  "0010011010010";
		Trees_din <= x"00054f08";
		wait for Clk_period;
		Addr <=  "0010011010011";
		Trees_din <= x"0a004104";
		wait for Clk_period;
		Addr <=  "0010011010100";
		Trees_din <= x"00361419";
		wait for Clk_period;
		Addr <=  "0010011010101";
		Trees_din <= x"ffa11419";
		wait for Clk_period;
		Addr <=  "0010011010110";
		Trees_din <= x"02072d04";
		wait for Clk_period;
		Addr <=  "0010011010111";
		Trees_din <= x"00e51419";
		wait for Clk_period;
		Addr <=  "0010011011000";
		Trees_din <= x"00081419";
		wait for Clk_period;
		Addr <=  "0010011011001";
		Trees_din <= x"04f99b0c";
		wait for Clk_period;
		Addr <=  "0010011011010";
		Trees_din <= x"03f81308";
		wait for Clk_period;
		Addr <=  "0010011011011";
		Trees_din <= x"0f001704";
		wait for Clk_period;
		Addr <=  "0010011011100";
		Trees_din <= x"013a1419";
		wait for Clk_period;
		Addr <=  "0010011011101";
		Trees_din <= x"00221419";
		wait for Clk_period;
		Addr <=  "0010011011110";
		Trees_din <= x"ff921419";
		wait for Clk_period;
		Addr <=  "0010011011111";
		Trees_din <= x"06fc2008";
		wait for Clk_period;
		Addr <=  "0010011100000";
		Trees_din <= x"0a004404";
		wait for Clk_period;
		Addr <=  "0010011100001";
		Trees_din <= x"006f1419";
		wait for Clk_period;
		Addr <=  "0010011100010";
		Trees_din <= x"ff911419";
		wait for Clk_period;
		Addr <=  "0010011100011";
		Trees_din <= x"0a005804";
		wait for Clk_period;
		Addr <=  "0010011100100";
		Trees_din <= x"ff711419";
		wait for Clk_period;
		Addr <=  "0010011100101";
		Trees_din <= x"fff31419";
		wait for Clk_period;
		Addr <=  "0010011100110";
		Trees_din <= x"0b009320";
		wait for Clk_period;
		Addr <=  "0010011100111";
		Trees_din <= x"0b007410";
		wait for Clk_period;
		Addr <=  "0010011101000";
		Trees_din <= x"0c00ae08";
		wait for Clk_period;
		Addr <=  "0010011101001";
		Trees_din <= x"03f89504";
		wait for Clk_period;
		Addr <=  "0010011101010";
		Trees_din <= x"00251419";
		wait for Clk_period;
		Addr <=  "0010011101011";
		Trees_din <= x"ffdb1419";
		wait for Clk_period;
		Addr <=  "0010011101100";
		Trees_din <= x"07f5b904";
		wait for Clk_period;
		Addr <=  "0010011101101";
		Trees_din <= x"ffaf1419";
		wait for Clk_period;
		Addr <=  "0010011101110";
		Trees_din <= x"006e1419";
		wait for Clk_period;
		Addr <=  "0010011101111";
		Trees_din <= x"03fa4608";
		wait for Clk_period;
		Addr <=  "0010011110000";
		Trees_din <= x"06fc9a04";
		wait for Clk_period;
		Addr <=  "0010011110001";
		Trees_din <= x"ff801419";
		wait for Clk_period;
		Addr <=  "0010011110010";
		Trees_din <= x"fffa1419";
		wait for Clk_period;
		Addr <=  "0010011110011";
		Trees_din <= x"0d014704";
		wait for Clk_period;
		Addr <=  "0010011110100";
		Trees_din <= x"00bf1419";
		wait for Clk_period;
		Addr <=  "0010011110101";
		Trees_din <= x"ffd91419";
		wait for Clk_period;
		Addr <=  "0010011110110";
		Trees_din <= x"1c028710";
		wait for Clk_period;
		Addr <=  "0010011110111";
		Trees_din <= x"04003a08";
		wait for Clk_period;
		Addr <=  "0010011111000";
		Trees_din <= x"2003fb04";
		wait for Clk_period;
		Addr <=  "0010011111001";
		Trees_din <= x"ff9f1419";
		wait for Clk_period;
		Addr <=  "0010011111010";
		Trees_din <= x"009d1419";
		wait for Clk_period;
		Addr <=  "0010011111011";
		Trees_din <= x"0c00d904";
		wait for Clk_period;
		Addr <=  "0010011111100";
		Trees_din <= x"ffce1419";
		wait for Clk_period;
		Addr <=  "0010011111101";
		Trees_din <= x"00651419";
		wait for Clk_period;
		Addr <=  "0010011111110";
		Trees_din <= x"0b009604";
		wait for Clk_period;
		Addr <=  "0010011111111";
		Trees_din <= x"00691419";
		wait for Clk_period;
		Addr <=  "0010100000000";
		Trees_din <= x"12008304";
		wait for Clk_period;
		Addr <=  "0010100000001";
		Trees_din <= x"ffd91419";
		wait for Clk_period;
		Addr <=  "0010100000010";
		Trees_din <= x"ff5a1419";
		wait for Clk_period;
		Addr <=  "0010100000011";
		Trees_din <= x"00178004";
		wait for Clk_period;
		Addr <=  "0010100000100";
		Trees_din <= x"00331419";
		wait for Clk_period;
		Addr <=  "0010100000101";
		Trees_din <= x"00981419";
		wait for Clk_period;
		Addr <=  "0010100000110";
		Trees_din <= x"0016b450";
		wait for Clk_period;
		Addr <=  "0010100000111";
		Trees_din <= x"00026914";
		wait for Clk_period;
		Addr <=  "0010100001000";
		Trees_din <= x"05f99f04";
		wait for Clk_period;
		Addr <=  "0010100001001";
		Trees_din <= x"ff7414c5";
		wait for Clk_period;
		Addr <=  "0010100001010";
		Trees_din <= x"05f9f504";
		wait for Clk_period;
		Addr <=  "0010100001011";
		Trees_din <= x"008e14c5";
		wait for Clk_period;
		Addr <=  "0010100001100";
		Trees_din <= x"04fad704";
		wait for Clk_period;
		Addr <=  "0010100001101";
		Trees_din <= x"ff7a14c5";
		wait for Clk_period;
		Addr <=  "0010100001110";
		Trees_din <= x"04fb6a04";
		wait for Clk_period;
		Addr <=  "0010100001111";
		Trees_din <= x"009f14c5";
		wait for Clk_period;
		Addr <=  "0010100010000";
		Trees_din <= x"ffd414c5";
		wait for Clk_period;
		Addr <=  "0010100010001";
		Trees_din <= x"06fb451c";
		wait for Clk_period;
		Addr <=  "0010100010010";
		Trees_din <= x"03f7de0c";
		wait for Clk_period;
		Addr <=  "0010100010011";
		Trees_din <= x"06faeb08";
		wait for Clk_period;
		Addr <=  "0010100010100";
		Trees_din <= x"1303ed04";
		wait for Clk_period;
		Addr <=  "0010100010101";
		Trees_din <= x"ff6214c5";
		wait for Clk_period;
		Addr <=  "0010100010110";
		Trees_din <= x"000a14c5";
		wait for Clk_period;
		Addr <=  "0010100010111";
		Trees_din <= x"005e14c5";
		wait for Clk_period;
		Addr <=  "0010100011000";
		Trees_din <= x"15004608";
		wait for Clk_period;
		Addr <=  "0010100011001";
		Trees_din <= x"13034904";
		wait for Clk_period;
		Addr <=  "0010100011010";
		Trees_din <= x"ffe714c5";
		wait for Clk_period;
		Addr <=  "0010100011011";
		Trees_din <= x"00c714c5";
		wait for Clk_period;
		Addr <=  "0010100011100";
		Trees_din <= x"0900c604";
		wait for Clk_period;
		Addr <=  "0010100011101";
		Trees_din <= x"ff8914c5";
		wait for Clk_period;
		Addr <=  "0010100011110";
		Trees_din <= x"fff714c5";
		wait for Clk_period;
		Addr <=  "0010100011111";
		Trees_din <= x"21000010";
		wait for Clk_period;
		Addr <=  "0010100100000";
		Trees_din <= x"0b007408";
		wait for Clk_period;
		Addr <=  "0010100100001";
		Trees_din <= x"12007c04";
		wait for Clk_period;
		Addr <=  "0010100100010";
		Trees_din <= x"000c14c5";
		wait for Clk_period;
		Addr <=  "0010100100011";
		Trees_din <= x"006614c5";
		wait for Clk_period;
		Addr <=  "0010100100100";
		Trees_din <= x"06fc8b04";
		wait for Clk_period;
		Addr <=  "0010100100101";
		Trees_din <= x"ff8214c5";
		wait for Clk_period;
		Addr <=  "0010100100110";
		Trees_din <= x"fffe14c5";
		wait for Clk_period;
		Addr <=  "0010100100111";
		Trees_din <= x"0b007d08";
		wait for Clk_period;
		Addr <=  "0010100101000";
		Trees_din <= x"07fe6604";
		wait for Clk_period;
		Addr <=  "0010100101001";
		Trees_din <= x"00b214c5";
		wait for Clk_period;
		Addr <=  "0010100101010";
		Trees_din <= x"ffd514c5";
		wait for Clk_period;
		Addr <=  "0010100101011";
		Trees_din <= x"17fa1104";
		wait for Clk_period;
		Addr <=  "0010100101100";
		Trees_din <= x"ffda14c5";
		wait for Clk_period;
		Addr <=  "0010100101101";
		Trees_din <= x"008814c5";
		wait for Clk_period;
		Addr <=  "0010100101110";
		Trees_din <= x"00178004";
		wait for Clk_period;
		Addr <=  "0010100101111";
		Trees_din <= x"003014c5";
		wait for Clk_period;
		Addr <=  "0010100110000";
		Trees_din <= x"009514c5";
		wait for Clk_period;
		Addr <=  "0010100110001";
		Trees_din <= x"0012e55c";
		wait for Clk_period;
		Addr <=  "0010100110010";
		Trees_din <= x"0006261c";
		wait for Clk_period;
		Addr <=  "0010100110011";
		Trees_din <= x"02083318";
		wait for Clk_period;
		Addr <=  "0010100110100";
		Trees_din <= x"0b008810";
		wait for Clk_period;
		Addr <=  "0010100110101";
		Trees_din <= x"010c3408";
		wait for Clk_period;
		Addr <=  "0010100110110";
		Trees_din <= x"0f000a04";
		wait for Clk_period;
		Addr <=  "0010100110111";
		Trees_din <= x"005015b1";
		wait for Clk_period;
		Addr <=  "0010100111000";
		Trees_din <= x"ffe215b1";
		wait for Clk_period;
		Addr <=  "0010100111001";
		Trees_din <= x"11024004";
		wait for Clk_period;
		Addr <=  "0010100111010";
		Trees_din <= x"ff7615b1";
		wait for Clk_period;
		Addr <=  "0010100111011";
		Trees_din <= x"002f15b1";
		wait for Clk_period;
		Addr <=  "0010100111100";
		Trees_din <= x"03028704";
		wait for Clk_period;
		Addr <=  "0010100111101";
		Trees_din <= x"ff7615b1";
		wait for Clk_period;
		Addr <=  "0010100111110";
		Trees_din <= x"001715b1";
		wait for Clk_period;
		Addr <=  "0010100111111";
		Trees_din <= x"ff7615b1";
		wait for Clk_period;
		Addr <=  "0010101000000";
		Trees_din <= x"0b008720";
		wait for Clk_period;
		Addr <=  "0010101000001";
		Trees_din <= x"03f69210";
		wait for Clk_period;
		Addr <=  "0010101000010";
		Trees_din <= x"07ff8f08";
		wait for Clk_period;
		Addr <=  "0010101000011";
		Trees_din <= x"03f66004";
		wait for Clk_period;
		Addr <=  "0010101000100";
		Trees_din <= x"000a15b1";
		wait for Clk_period;
		Addr <=  "0010101000101";
		Trees_din <= x"ff6615b1";
		wait for Clk_period;
		Addr <=  "0010101000110";
		Trees_din <= x"10003c04";
		wait for Clk_period;
		Addr <=  "0010101000111";
		Trees_din <= x"007015b1";
		wait for Clk_period;
		Addr <=  "0010101001000";
		Trees_din <= x"ff5915b1";
		wait for Clk_period;
		Addr <=  "0010101001001";
		Trees_din <= x"0b008408";
		wait for Clk_period;
		Addr <=  "0010101001010";
		Trees_din <= x"03f86004";
		wait for Clk_period;
		Addr <=  "0010101001011";
		Trees_din <= x"003315b1";
		wait for Clk_period;
		Addr <=  "0010101001100";
		Trees_din <= x"fffe15b1";
		wait for Clk_period;
		Addr <=  "0010101001101";
		Trees_din <= x"000f5404";
		wait for Clk_period;
		Addr <=  "0010101001110";
		Trees_din <= x"ff4d15b1";
		wait for Clk_period;
		Addr <=  "0010101001111";
		Trees_din <= x"006115b1";
		wait for Clk_period;
		Addr <=  "0010101010000";
		Trees_din <= x"03f50b10";
		wait for Clk_period;
		Addr <=  "0010101010001";
		Trees_din <= x"04003a08";
		wait for Clk_period;
		Addr <=  "0010101010010";
		Trees_din <= x"01106c04";
		wait for Clk_period;
		Addr <=  "0010101010011";
		Trees_din <= x"00f715b1";
		wait for Clk_period;
		Addr <=  "0010101010100";
		Trees_din <= x"fff415b1";
		wait for Clk_period;
		Addr <=  "0010101010101";
		Trees_din <= x"0b009004";
		wait for Clk_period;
		Addr <=  "0010101010110";
		Trees_din <= x"008c15b1";
		wait for Clk_period;
		Addr <=  "0010101010111";
		Trees_din <= x"ff8215b1";
		wait for Clk_period;
		Addr <=  "0010101011000";
		Trees_din <= x"1101b808";
		wait for Clk_period;
		Addr <=  "0010101011001";
		Trees_din <= x"11018504";
		wait for Clk_period;
		Addr <=  "0010101011010";
		Trees_din <= x"001c15b1";
		wait for Clk_period;
		Addr <=  "0010101011011";
		Trees_din <= x"00c615b1";
		wait for Clk_period;
		Addr <=  "0010101011100";
		Trees_din <= x"15003704";
		wait for Clk_period;
		Addr <=  "0010101011101";
		Trees_din <= x"ff7815b1";
		wait for Clk_period;
		Addr <=  "0010101011110";
		Trees_din <= x"001015b1";
		wait for Clk_period;
		Addr <=  "0010101011111";
		Trees_din <= x"0c00a804";
		wait for Clk_period;
		Addr <=  "0010101100000";
		Trees_din <= x"009115b1";
		wait for Clk_period;
		Addr <=  "0010101100001";
		Trees_din <= x"0c00ad08";
		wait for Clk_period;
		Addr <=  "0010101100010";
		Trees_din <= x"0401f404";
		wait for Clk_period;
		Addr <=  "0010101100011";
		Trees_din <= x"ff5215b1";
		wait for Clk_period;
		Addr <=  "0010101100100";
		Trees_din <= x"001815b1";
		wait for Clk_period;
		Addr <=  "0010101100101";
		Trees_din <= x"1e02870c";
		wait for Clk_period;
		Addr <=  "0010101100110";
		Trees_din <= x"01130b08";
		wait for Clk_period;
		Addr <=  "0010101100111";
		Trees_din <= x"0b00a204";
		wait for Clk_period;
		Addr <=  "0010101101000";
		Trees_din <= x"008c15b1";
		wait for Clk_period;
		Addr <=  "0010101101001";
		Trees_din <= x"001515b1";
		wait for Clk_period;
		Addr <=  "0010101101010";
		Trees_din <= x"000e15b1";
		wait for Clk_period;
		Addr <=  "0010101101011";
		Trees_din <= x"ffc115b1";
		wait for Clk_period;
		Addr <=  "0010101101100";
		Trees_din <= x"0016b430";
		wait for Clk_period;
		Addr <=  "0010101101101";
		Trees_din <= x"00fef408";
		wait for Clk_period;
		Addr <=  "0010101101110";
		Trees_din <= x"04fdb904";
		wait for Clk_period;
		Addr <=  "0010101101111";
		Trees_din <= x"ff7c1615";
		wait for Clk_period;
		Addr <=  "0010101110000";
		Trees_din <= x"00191615";
		wait for Clk_period;
		Addr <=  "0010101110001";
		Trees_din <= x"01f76408";
		wait for Clk_period;
		Addr <=  "0010101110010";
		Trees_din <= x"0900b304";
		wait for Clk_period;
		Addr <=  "0010101110011";
		Trees_din <= x"00181615";
		wait for Clk_period;
		Addr <=  "0010101110100";
		Trees_din <= x"ff641615";
		wait for Clk_period;
		Addr <=  "0010101110101";
		Trees_din <= x"01046510";
		wait for Clk_period;
		Addr <=  "0010101110110";
		Trees_din <= x"0601f908";
		wait for Clk_period;
		Addr <=  "0010101110111";
		Trees_din <= x"0008df04";
		wait for Clk_period;
		Addr <=  "0010101111000";
		Trees_din <= x"ff8c1615";
		wait for Clk_period;
		Addr <=  "0010101111001";
		Trees_din <= x"001a1615";
		wait for Clk_period;
		Addr <=  "0010101111010";
		Trees_din <= x"0a004304";
		wait for Clk_period;
		Addr <=  "0010101111011";
		Trees_din <= x"00a61615";
		wait for Clk_period;
		Addr <=  "0010101111100";
		Trees_din <= x"fffd1615";
		wait for Clk_period;
		Addr <=  "0010101111101";
		Trees_din <= x"020a3108";
		wait for Clk_period;
		Addr <=  "0010101111110";
		Trees_din <= x"1b073c04";
		wait for Clk_period;
		Addr <=  "0010101111111";
		Trees_din <= x"00091615";
		wait for Clk_period;
		Addr <=  "0010110000000";
		Trees_din <= x"008c1615";
		wait for Clk_period;
		Addr <=  "0010110000001";
		Trees_din <= x"03f4a504";
		wait for Clk_period;
		Addr <=  "0010110000010";
		Trees_din <= x"00491615";
		wait for Clk_period;
		Addr <=  "0010110000011";
		Trees_din <= x"ffa01615";
		wait for Clk_period;
		Addr <=  "0010110000100";
		Trees_din <= x"00851615";
		wait for Clk_period;
		Addr <=  "0010110000101";
		Trees_din <= x"00178060";
		wait for Clk_period;
		Addr <=  "0010110000110";
		Trees_din <= x"0003b420";
		wait for Clk_period;
		Addr <=  "0010110000111";
		Trees_din <= x"02003c0c";
		wait for Clk_period;
		Addr <=  "0010110001000";
		Trees_din <= x"1afc5408";
		wait for Clk_period;
		Addr <=  "0010110001001";
		Trees_din <= x"1100e504";
		wait for Clk_period;
		Addr <=  "0010110001010";
		Trees_din <= x"00c716d9";
		wait for Clk_period;
		Addr <=  "0010110001011";
		Trees_din <= x"000816d9";
		wait for Clk_period;
		Addr <=  "0010110001100";
		Trees_din <= x"ff9c16d9";
		wait for Clk_period;
		Addr <=  "0010110001101";
		Trees_din <= x"0e003908";
		wait for Clk_period;
		Addr <=  "0010110001110";
		Trees_din <= x"01fc8c04";
		wait for Clk_period;
		Addr <=  "0010110001111";
		Trees_din <= x"001016d9";
		wait for Clk_period;
		Addr <=  "0010110010000";
		Trees_din <= x"ff6e16d9";
		wait for Clk_period;
		Addr <=  "0010110010001";
		Trees_din <= x"0108e508";
		wait for Clk_period;
		Addr <=  "0010110010010";
		Trees_din <= x"0f000904";
		wait for Clk_period;
		Addr <=  "0010110010011";
		Trees_din <= x"007916d9";
		wait for Clk_period;
		Addr <=  "0010110010100";
		Trees_din <= x"ffa116d9";
		wait for Clk_period;
		Addr <=  "0010110010101";
		Trees_din <= x"ff8b16d9";
		wait for Clk_period;
		Addr <=  "0010110010110";
		Trees_din <= x"04ff0d20";
		wait for Clk_period;
		Addr <=  "0010110010111";
		Trees_din <= x"06fcca10";
		wait for Clk_period;
		Addr <=  "0010110011000";
		Trees_din <= x"19001608";
		wait for Clk_period;
		Addr <=  "0010110011001";
		Trees_din <= x"15004604";
		wait for Clk_period;
		Addr <=  "0010110011010";
		Trees_din <= x"008e16d9";
		wait for Clk_period;
		Addr <=  "0010110011011";
		Trees_din <= x"ffd216d9";
		wait for Clk_period;
		Addr <=  "0010110011100";
		Trees_din <= x"1b028204";
		wait for Clk_period;
		Addr <=  "0010110011101";
		Trees_din <= x"ff6216d9";
		wait for Clk_period;
		Addr <=  "0010110011110";
		Trees_din <= x"ffe616d9";
		wait for Clk_period;
		Addr <=  "0010110011111";
		Trees_din <= x"07fe7408";
		wait for Clk_period;
		Addr <=  "0010110100000";
		Trees_din <= x"010cb704";
		wait for Clk_period;
		Addr <=  "0010110100001";
		Trees_din <= x"004d16d9";
		wait for Clk_period;
		Addr <=  "0010110100010";
		Trees_din <= x"fffd16d9";
		wait for Clk_period;
		Addr <=  "0010110100011";
		Trees_din <= x"15003104";
		wait for Clk_period;
		Addr <=  "0010110100100";
		Trees_din <= x"006916d9";
		wait for Clk_period;
		Addr <=  "0010110100101";
		Trees_din <= x"ffd616d9";
		wait for Clk_period;
		Addr <=  "0010110100110";
		Trees_din <= x"20040010";
		wait for Clk_period;
		Addr <=  "0010110100111";
		Trees_din <= x"14040008";
		wait for Clk_period;
		Addr <=  "0010110101000";
		Trees_din <= x"14040004";
		wait for Clk_period;
		Addr <=  "0010110101001";
		Trees_din <= x"002816d9";
		wait for Clk_period;
		Addr <=  "0010110101010";
		Trees_din <= x"00de16d9";
		wait for Clk_period;
		Addr <=  "0010110101011";
		Trees_din <= x"000f7304";
		wait for Clk_period;
		Addr <=  "0010110101100";
		Trees_din <= x"ff4916d9";
		wait for Clk_period;
		Addr <=  "0010110101101";
		Trees_din <= x"003116d9";
		wait for Clk_period;
		Addr <=  "0010110101110";
		Trees_din <= x"01083708";
		wait for Clk_period;
		Addr <=  "0010110101111";
		Trees_din <= x"03f9af04";
		wait for Clk_period;
		Addr <=  "0010110110000";
		Trees_din <= x"fffc16d9";
		wait for Clk_period;
		Addr <=  "0010110110001";
		Trees_din <= x"008316d9";
		wait for Clk_period;
		Addr <=  "0010110110010";
		Trees_din <= x"05f68e04";
		wait for Clk_period;
		Addr <=  "0010110110011";
		Trees_din <= x"fff616d9";
		wait for Clk_period;
		Addr <=  "0010110110100";
		Trees_din <= x"ff7e16d9";
		wait for Clk_period;
		Addr <=  "0010110110101";
		Trees_din <= x"008916d9";
		wait for Clk_period;
		Addr <=  "0010110110110";
		Trees_din <= x"0016b460";
		wait for Clk_period;
		Addr <=  "0010110110111";
		Trees_din <= x"0405f140";
		wait for Clk_period;
		Addr <=  "0010110111000";
		Trees_din <= x"0009b220";
		wait for Clk_period;
		Addr <=  "0010110111001";
		Trees_din <= x"0c00c310";
		wait for Clk_period;
		Addr <=  "0010110111010";
		Trees_din <= x"08003808";
		wait for Clk_period;
		Addr <=  "0010110111011";
		Trees_din <= x"04f95a04";
		wait for Clk_period;
		Addr <=  "0010110111100";
		Trees_din <= x"007a179d";
		wait for Clk_period;
		Addr <=  "0010110111101";
		Trees_din <= x"ff84179d";
		wait for Clk_period;
		Addr <=  "0010110111110";
		Trees_din <= x"03f75704";
		wait for Clk_period;
		Addr <=  "0010110111111";
		Trees_din <= x"ffaa179d";
		wait for Clk_period;
		Addr <=  "0010111000000";
		Trees_din <= x"000a179d";
		wait for Clk_period;
		Addr <=  "0010111000001";
		Trees_din <= x"0c00dc08";
		wait for Clk_period;
		Addr <=  "0010111000010";
		Trees_din <= x"03f84004";
		wait for Clk_period;
		Addr <=  "0010111000011";
		Trees_din <= x"00d3179d";
		wait for Clk_period;
		Addr <=  "0010111000100";
		Trees_din <= x"000c179d";
		wait for Clk_period;
		Addr <=  "0010111000101";
		Trees_din <= x"00081904";
		wait for Clk_period;
		Addr <=  "0010111000110";
		Trees_din <= x"ff66179d";
		wait for Clk_period;
		Addr <=  "0010111000111";
		Trees_din <= x"0038179d";
		wait for Clk_period;
		Addr <=  "0010111001000";
		Trees_din <= x"0c009e10";
		wait for Clk_period;
		Addr <=  "0010111001001";
		Trees_din <= x"06003508";
		wait for Clk_period;
		Addr <=  "0010111001010";
		Trees_din <= x"16009604";
		wait for Clk_period;
		Addr <=  "0010111001011";
		Trees_din <= x"0058179d";
		wait for Clk_period;
		Addr <=  "0010111001100";
		Trees_din <= x"ffe1179d";
		wait for Clk_period;
		Addr <=  "0010111001101";
		Trees_din <= x"0602d004";
		wait for Clk_period;
		Addr <=  "0010111001110";
		Trees_din <= x"ffd4179d";
		wait for Clk_period;
		Addr <=  "0010111001111";
		Trees_din <= x"0056179d";
		wait for Clk_period;
		Addr <=  "0010111010000";
		Trees_din <= x"0c00a008";
		wait for Clk_period;
		Addr <=  "0010111010001";
		Trees_din <= x"08004704";
		wait for Clk_period;
		Addr <=  "0010111010010";
		Trees_din <= x"ff5d179d";
		wait for Clk_period;
		Addr <=  "0010111010011";
		Trees_din <= x"0092179d";
		wait for Clk_period;
		Addr <=  "0010111010100";
		Trees_din <= x"0600c904";
		wait for Clk_period;
		Addr <=  "0010111010101";
		Trees_din <= x"0000179d";
		wait for Clk_period;
		Addr <=  "0010111010110";
		Trees_din <= x"0037179d";
		wait for Clk_period;
		Addr <=  "0010111010111";
		Trees_din <= x"03fa4618";
		wait for Clk_period;
		Addr <=  "0010111011000";
		Trees_din <= x"00114810";
		wait for Clk_period;
		Addr <=  "0010111011001";
		Trees_din <= x"0b008508";
		wait for Clk_period;
		Addr <=  "0010111011010";
		Trees_din <= x"0f005804";
		wait for Clk_period;
		Addr <=  "0010111011011";
		Trees_din <= x"ff4a179d";
		wait for Clk_period;
		Addr <=  "0010111011100";
		Trees_din <= x"0020179d";
		wait for Clk_period;
		Addr <=  "0010111011101";
		Trees_din <= x"07f75e04";
		wait for Clk_period;
		Addr <=  "0010111011110";
		Trees_din <= x"ff9a179d";
		wait for Clk_period;
		Addr <=  "0010111011111";
		Trees_din <= x"0072179d";
		wait for Clk_period;
		Addr <=  "0010111100000";
		Trees_din <= x"10003304";
		wait for Clk_period;
		Addr <=  "0010111100001";
		Trees_din <= x"ffa4179d";
		wait for Clk_period;
		Addr <=  "0010111100010";
		Trees_din <= x"0078179d";
		wait for Clk_period;
		Addr <=  "0010111100011";
		Trees_din <= x"14040004";
		wait for Clk_period;
		Addr <=  "0010111100100";
		Trees_din <= x"0016179d";
		wait for Clk_period;
		Addr <=  "0010111100101";
		Trees_din <= x"0078179d";
		wait for Clk_period;
		Addr <=  "0010111100110";
		Trees_din <= x"007c179d";
		wait for Clk_period;
		Addr <=  "0010111100111";
		Trees_din <= x"000fee70";
		wait for Clk_period;
		Addr <=  "0010111101000";
		Trees_din <= x"0a004734";
		wait for Clk_period;
		Addr <=  "0010111101001";
		Trees_din <= x"0900b518";
		wait for Clk_period;
		Addr <=  "0010111101010";
		Trees_din <= x"02093410";
		wait for Clk_period;
		Addr <=  "0010111101011";
		Trees_din <= x"010f2f08";
		wait for Clk_period;
		Addr <=  "0010111101100";
		Trees_din <= x"1b027304";
		wait for Clk_period;
		Addr <=  "0010111101101";
		Trees_din <= x"004a1911";
		wait for Clk_period;
		Addr <=  "0010111101110";
		Trees_din <= x"00c71911";
		wait for Clk_period;
		Addr <=  "0010111101111";
		Trees_din <= x"06010204";
		wait for Clk_period;
		Addr <=  "0010111110000";
		Trees_din <= x"ff911911";
		wait for Clk_period;
		Addr <=  "0010111110001";
		Trees_din <= x"00771911";
		wait for Clk_period;
		Addr <=  "0010111110010";
		Trees_din <= x"07f85a04";
		wait for Clk_period;
		Addr <=  "0010111110011";
		Trees_din <= x"ffdd1911";
		wait for Clk_period;
		Addr <=  "0010111110100";
		Trees_din <= x"ff771911";
		wait for Clk_period;
		Addr <=  "0010111110101";
		Trees_din <= x"0900ba0c";
		wait for Clk_period;
		Addr <=  "0010111110110";
		Trees_din <= x"06fc5f04";
		wait for Clk_period;
		Addr <=  "0010111110111";
		Trees_din <= x"00861911";
		wait for Clk_period;
		Addr <=  "0010111111000";
		Trees_din <= x"000ca304";
		wait for Clk_period;
		Addr <=  "0010111111001";
		Trees_din <= x"ff531911";
		wait for Clk_period;
		Addr <=  "0010111111010";
		Trees_din <= x"000d1911";
		wait for Clk_period;
		Addr <=  "0010111111011";
		Trees_din <= x"18005208";
		wait for Clk_period;
		Addr <=  "0010111111100";
		Trees_din <= x"11018b04";
		wait for Clk_period;
		Addr <=  "0010111111101";
		Trees_din <= x"00171911";
		wait for Clk_period;
		Addr <=  "0010111111110";
		Trees_din <= x"00ba1911";
		wait for Clk_period;
		Addr <=  "0010111111111";
		Trees_din <= x"1403e704";
		wait for Clk_period;
		Addr <=  "0011000000000";
		Trees_din <= x"000f1911";
		wait for Clk_period;
		Addr <=  "0011000000001";
		Trees_din <= x"ffca1911";
		wait for Clk_period;
		Addr <=  "0011000000010";
		Trees_din <= x"0a004f20";
		wait for Clk_period;
		Addr <=  "0011000000011";
		Trees_din <= x"02033910";
		wait for Clk_period;
		Addr <=  "0011000000100";
		Trees_din <= x"06febc08";
		wait for Clk_period;
		Addr <=  "0011000000101";
		Trees_din <= x"10004a04";
		wait for Clk_period;
		Addr <=  "0011000000110";
		Trees_din <= x"00ce1911";
		wait for Clk_period;
		Addr <=  "0011000000111";
		Trees_din <= x"fffd1911";
		wait for Clk_period;
		Addr <=  "0011000001000";
		Trees_din <= x"06013d04";
		wait for Clk_period;
		Addr <=  "0011000001001";
		Trees_din <= x"ff641911";
		wait for Clk_period;
		Addr <=  "0011000001010";
		Trees_din <= x"004a1911";
		wait for Clk_period;
		Addr <=  "0011000001011";
		Trees_din <= x"000b5708";
		wait for Clk_period;
		Addr <=  "0011000001100";
		Trees_din <= x"0c00a004";
		wait for Clk_period;
		Addr <=  "0011000001101";
		Trees_din <= x"ffe91911";
		wait for Clk_period;
		Addr <=  "0011000001110";
		Trees_din <= x"ff791911";
		wait for Clk_period;
		Addr <=  "0011000001111";
		Trees_din <= x"15003e04";
		wait for Clk_period;
		Addr <=  "0011000010000";
		Trees_din <= x"003d1911";
		wait for Clk_period;
		Addr <=  "0011000010001";
		Trees_din <= x"ffbe1911";
		wait for Clk_period;
		Addr <=  "0011000010010";
		Trees_din <= x"0104b10c";
		wait for Clk_period;
		Addr <=  "0011000010011";
		Trees_din <= x"01faca04";
		wait for Clk_period;
		Addr <=  "0011000010100";
		Trees_din <= x"00481911";
		wait for Clk_period;
		Addr <=  "0011000010101";
		Trees_din <= x"000bb504";
		wait for Clk_period;
		Addr <=  "0011000010110";
		Trees_din <= x"ff461911";
		wait for Clk_period;
		Addr <=  "0011000010111";
		Trees_din <= x"ffe21911";
		wait for Clk_period;
		Addr <=  "0011000011000";
		Trees_din <= x"15004508";
		wait for Clk_period;
		Addr <=  "0011000011001";
		Trees_din <= x"12008504";
		wait for Clk_period;
		Addr <=  "0011000011010";
		Trees_din <= x"00aa1911";
		wait for Clk_period;
		Addr <=  "0011000011011";
		Trees_din <= x"00151911";
		wait for Clk_period;
		Addr <=  "0011000011100";
		Trees_din <= x"17fff904";
		wait for Clk_period;
		Addr <=  "0011000011101";
		Trees_din <= x"ffd51911";
		wait for Clk_period;
		Addr <=  "0011000011110";
		Trees_din <= x"00991911";
		wait for Clk_period;
		Addr <=  "0011000011111";
		Trees_din <= x"0a004330";
		wait for Clk_period;
		Addr <=  "0011000100000";
		Trees_din <= x"0a003f14";
		wait for Clk_period;
		Addr <=  "0011000100001";
		Trees_din <= x"0d000404";
		wait for Clk_period;
		Addr <=  "0011000100010";
		Trees_din <= x"ff9e1911";
		wait for Clk_period;
		Addr <=  "0011000100011";
		Trees_din <= x"0900bb08";
		wait for Clk_period;
		Addr <=  "0011000100100";
		Trees_din <= x"11018904";
		wait for Clk_period;
		Addr <=  "0011000100101";
		Trees_din <= x"ff881911";
		wait for Clk_period;
		Addr <=  "0011000100110";
		Trees_din <= x"003e1911";
		wait for Clk_period;
		Addr <=  "0011000100111";
		Trees_din <= x"05f75104";
		wait for Clk_period;
		Addr <=  "0011000101000";
		Trees_din <= x"008b1911";
		wait for Clk_period;
		Addr <=  "0011000101001";
		Trees_din <= x"ffc41911";
		wait for Clk_period;
		Addr <=  "0011000101010";
		Trees_din <= x"00110d0c";
		wait for Clk_period;
		Addr <=  "0011000101011";
		Trees_din <= x"08004508";
		wait for Clk_period;
		Addr <=  "0011000101100";
		Trees_din <= x"08003c04";
		wait for Clk_period;
		Addr <=  "0011000101101";
		Trees_din <= x"fff21911";
		wait for Clk_period;
		Addr <=  "0011000101110";
		Trees_din <= x"ff011911";
		wait for Clk_period;
		Addr <=  "0011000101111";
		Trees_din <= x"00571911";
		wait for Clk_period;
		Addr <=  "0011000110000";
		Trees_din <= x"010dac08";
		wait for Clk_period;
		Addr <=  "0011000110001";
		Trees_din <= x"03f70b04";
		wait for Clk_period;
		Addr <=  "0011000110010";
		Trees_din <= x"00871911";
		wait for Clk_period;
		Addr <=  "0011000110011";
		Trees_din <= x"ffc91911";
		wait for Clk_period;
		Addr <=  "0011000110100";
		Trees_din <= x"1302eb04";
		wait for Clk_period;
		Addr <=  "0011000110101";
		Trees_din <= x"00161911";
		wait for Clk_period;
		Addr <=  "0011000110110";
		Trees_din <= x"ff861911";
		wait for Clk_period;
		Addr <=  "0011000110111";
		Trees_din <= x"18031c14";
		wait for Clk_period;
		Addr <=  "0011000111000";
		Trees_din <= x"11016a0c";
		wait for Clk_period;
		Addr <=  "0011000111001";
		Trees_din <= x"11014808";
		wait for Clk_period;
		Addr <=  "0011000111010";
		Trees_din <= x"08003704";
		wait for Clk_period;
		Addr <=  "0011000111011";
		Trees_din <= x"00001911";
		wait for Clk_period;
		Addr <=  "0011000111100";
		Trees_din <= x"00691911";
		wait for Clk_period;
		Addr <=  "0011000111101";
		Trees_din <= x"ff8b1911";
		wait for Clk_period;
		Addr <=  "0011000111110";
		Trees_din <= x"01110304";
		wait for Clk_period;
		Addr <=  "0011000111111";
		Trees_din <= x"009c1911";
		wait for Clk_period;
		Addr <=  "0011001000000";
		Trees_din <= x"ffec1911";
		wait for Clk_period;
		Addr <=  "0011001000001";
		Trees_din <= x"10003a04";
		wait for Clk_period;
		Addr <=  "0011001000010";
		Trees_din <= x"ff5a1911";
		wait for Clk_period;
		Addr <=  "0011001000011";
		Trees_din <= x"00021911";
		wait for Clk_period;
		Addr <=  "0011001000100";
		Trees_din <= x"00178044";
		wait for Clk_period;
		Addr <=  "0011001000101";
		Trees_din <= x"13008808";
		wait for Clk_period;
		Addr <=  "0011001000110";
		Trees_din <= x"0206c404";
		wait for Clk_period;
		Addr <=  "0011001000111";
		Trees_din <= x"fffc199d";
		wait for Clk_period;
		Addr <=  "0011001001000";
		Trees_din <= x"00bb199d";
		wait for Clk_period;
		Addr <=  "0011001001001";
		Trees_din <= x"0007e61c";
		wait for Clk_period;
		Addr <=  "0011001001010";
		Trees_din <= x"0900ad0c";
		wait for Clk_period;
		Addr <=  "0011001001011";
		Trees_din <= x"1403fa08";
		wait for Clk_period;
		Addr <=  "0011001001100";
		Trees_din <= x"05f6cc04";
		wait for Clk_period;
		Addr <=  "0011001001101";
		Trees_din <= x"ff71199d";
		wait for Clk_period;
		Addr <=  "0011001001110";
		Trees_din <= x"0019199d";
		wait for Clk_period;
		Addr <=  "0011001001111";
		Trees_din <= x"ff69199d";
		wait for Clk_period;
		Addr <=  "0011001010000";
		Trees_din <= x"0e003208";
		wait for Clk_period;
		Addr <=  "0011001010001";
		Trees_din <= x"0e002b04";
		wait for Clk_period;
		Addr <=  "0011001010010";
		Trees_din <= x"000e199d";
		wait for Clk_period;
		Addr <=  "0011001010011";
		Trees_din <= x"ff7a199d";
		wait for Clk_period;
		Addr <=  "0011001010100";
		Trees_din <= x"15004904";
		wait for Clk_period;
		Addr <=  "0011001010101";
		Trees_din <= x"0055199d";
		wait for Clk_period;
		Addr <=  "0011001010110";
		Trees_din <= x"ffc1199d";
		wait for Clk_period;
		Addr <=  "0011001010111";
		Trees_din <= x"00083c10";
		wait for Clk_period;
		Addr <=  "0011001011000";
		Trees_din <= x"03f7a908";
		wait for Clk_period;
		Addr <=  "0011001011001";
		Trees_din <= x"0f000404";
		wait for Clk_period;
		Addr <=  "0011001011010";
		Trees_din <= x"fffc199d";
		wait for Clk_period;
		Addr <=  "0011001011011";
		Trees_din <= x"ff65199d";
		wait for Clk_period;
		Addr <=  "0011001011100";
		Trees_din <= x"0f004b04";
		wait for Clk_period;
		Addr <=  "0011001011101";
		Trees_din <= x"00c2199d";
		wait for Clk_period;
		Addr <=  "0011001011110";
		Trees_din <= x"ffc4199d";
		wait for Clk_period;
		Addr <=  "0011001011111";
		Trees_din <= x"11000008";
		wait for Clk_period;
		Addr <=  "0011001100000";
		Trees_din <= x"12006704";
		wait for Clk_period;
		Addr <=  "0011001100001";
		Trees_din <= x"ffbe199d";
		wait for Clk_period;
		Addr <=  "0011001100010";
		Trees_din <= x"00b1199d";
		wait for Clk_period;
		Addr <=  "0011001100011";
		Trees_din <= x"01044d04";
		wait for Clk_period;
		Addr <=  "0011001100100";
		Trees_din <= x"002f199d";
		wait for Clk_period;
		Addr <=  "0011001100101";
		Trees_din <= x"ffff199d";
		wait for Clk_period;
		Addr <=  "0011001100110";
		Trees_din <= x"007f199d";
		wait for Clk_period;
		Addr <=  "0011001100111";
		Trees_din <= x"0003b428";
		wait for Clk_period;
		Addr <=  "0011001101000";
		Trees_din <= x"0108e520";
		wait for Clk_period;
		Addr <=  "0011001101001";
		Trees_din <= x"19000414";
		wait for Clk_period;
		Addr <=  "0011001101010";
		Trees_din <= x"0c008508";
		wait for Clk_period;
		Addr <=  "0011001101011";
		Trees_din <= x"0d013504";
		wait for Clk_period;
		Addr <=  "0011001101100";
		Trees_din <= x"ffee1aa9";
		wait for Clk_period;
		Addr <=  "0011001101101";
		Trees_din <= x"00831aa9";
		wait for Clk_period;
		Addr <=  "0011001101110";
		Trees_din <= x"0900b408";
		wait for Clk_period;
		Addr <=  "0011001101111";
		Trees_din <= x"0a004304";
		wait for Clk_period;
		Addr <=  "0011001110000";
		Trees_din <= x"007e1aa9";
		wait for Clk_period;
		Addr <=  "0011001110001";
		Trees_din <= x"ff8b1aa9";
		wait for Clk_period;
		Addr <=  "0011001110010";
		Trees_din <= x"ff7e1aa9";
		wait for Clk_period;
		Addr <=  "0011001110011";
		Trees_din <= x"17f8c208";
		wait for Clk_period;
		Addr <=  "0011001110100";
		Trees_din <= x"12007904";
		wait for Clk_period;
		Addr <=  "0011001110101";
		Trees_din <= x"00b91aa9";
		wait for Clk_period;
		Addr <=  "0011001110110";
		Trees_din <= x"002f1aa9";
		wait for Clk_period;
		Addr <=  "0011001110111";
		Trees_din <= x"ffa41aa9";
		wait for Clk_period;
		Addr <=  "0011001111000";
		Trees_din <= x"00036a04";
		wait for Clk_period;
		Addr <=  "0011001111001";
		Trees_din <= x"ff761aa9";
		wait for Clk_period;
		Addr <=  "0011001111010";
		Trees_din <= x"00111aa9";
		wait for Clk_period;
		Addr <=  "0011001111011";
		Trees_din <= x"04fe0c38";
		wait for Clk_period;
		Addr <=  "0011001111100";
		Trees_din <= x"1900051c";
		wait for Clk_period;
		Addr <=  "0011001111101";
		Trees_din <= x"0d02a210";
		wait for Clk_period;
		Addr <=  "0011001111110";
		Trees_din <= x"07fade08";
		wait for Clk_period;
		Addr <=  "0011001111111";
		Trees_din <= x"17f81a04";
		wait for Clk_period;
		Addr <=  "0011010000000";
		Trees_din <= x"00ab1aa9";
		wait for Clk_period;
		Addr <=  "0011010000001";
		Trees_din <= x"ff7d1aa9";
		wait for Clk_period;
		Addr <=  "0011010000010";
		Trees_din <= x"07fbfd04";
		wait for Clk_period;
		Addr <=  "0011010000011";
		Trees_din <= x"ff981aa9";
		wait for Clk_period;
		Addr <=  "0011010000100";
		Trees_din <= x"001e1aa9";
		wait for Clk_period;
		Addr <=  "0011010000101";
		Trees_din <= x"11020e08";
		wait for Clk_period;
		Addr <=  "0011010000110";
		Trees_din <= x"010d1604";
		wait for Clk_period;
		Addr <=  "0011010000111";
		Trees_din <= x"006a1aa9";
		wait for Clk_period;
		Addr <=  "0011010001000";
		Trees_din <= x"ffa31aa9";
		wait for Clk_period;
		Addr <=  "0011010001001";
		Trees_din <= x"01211aa9";
		wait for Clk_period;
		Addr <=  "0011010001010";
		Trees_din <= x"0f00880c";
		wait for Clk_period;
		Addr <=  "0011010001011";
		Trees_din <= x"03f5ec04";
		wait for Clk_period;
		Addr <=  "0011010001100";
		Trees_din <= x"00711aa9";
		wait for Clk_period;
		Addr <=  "0011010001101";
		Trees_din <= x"0a003c04";
		wait for Clk_period;
		Addr <=  "0011010001110";
		Trees_din <= x"00041aa9";
		wait for Clk_period;
		Addr <=  "0011010001111";
		Trees_din <= x"ff611aa9";
		wait for Clk_period;
		Addr <=  "0011010010000";
		Trees_din <= x"1b028608";
		wait for Clk_period;
		Addr <=  "0011010010001";
		Trees_din <= x"19000704";
		wait for Clk_period;
		Addr <=  "0011010010010";
		Trees_din <= x"ff721aa9";
		wait for Clk_period;
		Addr <=  "0011010010011";
		Trees_din <= x"007b1aa9";
		wait for Clk_period;
		Addr <=  "0011010010100";
		Trees_din <= x"04fd7504";
		wait for Clk_period;
		Addr <=  "0011010010101";
		Trees_din <= x"ff751aa9";
		wait for Clk_period;
		Addr <=  "0011010010110";
		Trees_din <= x"005a1aa9";
		wait for Clk_period;
		Addr <=  "0011010010111";
		Trees_din <= x"00066e0c";
		wait for Clk_period;
		Addr <=  "0011010011000";
		Trees_din <= x"1f023c04";
		wait for Clk_period;
		Addr <=  "0011010011001";
		Trees_din <= x"00121aa9";
		wait for Clk_period;
		Addr <=  "0011010011010";
		Trees_din <= x"0a005904";
		wait for Clk_period;
		Addr <=  "0011010011011";
		Trees_din <= x"ff731aa9";
		wait for Clk_period;
		Addr <=  "0011010011100";
		Trees_din <= x"000a1aa9";
		wait for Clk_period;
		Addr <=  "0011010011101";
		Trees_din <= x"0108640c";
		wait for Clk_period;
		Addr <=  "0011010011110";
		Trees_din <= x"04fe4a04";
		wait for Clk_period;
		Addr <=  "0011010011111";
		Trees_din <= x"ff581aa9";
		wait for Clk_period;
		Addr <=  "0011010100000";
		Trees_din <= x"1f028804";
		wait for Clk_period;
		Addr <=  "0011010100001";
		Trees_din <= x"002b1aa9";
		wait for Clk_period;
		Addr <=  "0011010100010";
		Trees_din <= x"ff811aa9";
		wait for Clk_period;
		Addr <=  "0011010100011";
		Trees_din <= x"0208a608";
		wait for Clk_period;
		Addr <=  "0011010100100";
		Trees_din <= x"05f69804";
		wait for Clk_period;
		Addr <=  "0011010100101";
		Trees_din <= x"000b1aa9";
		wait for Clk_period;
		Addr <=  "0011010100110";
		Trees_din <= x"ffbc1aa9";
		wait for Clk_period;
		Addr <=  "0011010100111";
		Trees_din <= x"06001504";
		wait for Clk_period;
		Addr <=  "0011010101000";
		Trees_din <= x"ffff1aa9";
		wait for Clk_period;
		Addr <=  "0011010101001";
		Trees_din <= x"ff751aa9";
		wait for Clk_period;
		Addr <=  "0011010101010";
		Trees_din <= x"0011e860";
		wait for Clk_period;
		Addr <=  "0011010101011";
		Trees_din <= x"07f5b924";
		wait for Clk_period;
		Addr <=  "0011010101100";
		Trees_din <= x"10004a14";
		wait for Clk_period;
		Addr <=  "0011010101101";
		Trees_din <= x"15003608";
		wait for Clk_period;
		Addr <=  "0011010101110";
		Trees_din <= x"08004004";
		wait for Clk_period;
		Addr <=  "0011010101111";
		Trees_din <= x"ffdf1bbd";
		wait for Clk_period;
		Addr <=  "0011010110000";
		Trees_din <= x"005f1bbd";
		wait for Clk_period;
		Addr <=  "0011010110001";
		Trees_din <= x"04ffbc04";
		wait for Clk_period;
		Addr <=  "0011010110010";
		Trees_din <= x"00021bbd";
		wait for Clk_period;
		Addr <=  "0011010110011";
		Trees_din <= x"1b025804";
		wait for Clk_period;
		Addr <=  "0011010110100";
		Trees_din <= x"00011bbd";
		wait for Clk_period;
		Addr <=  "0011010110101";
		Trees_din <= x"ff481bbd";
		wait for Clk_period;
		Addr <=  "0011010110110";
		Trees_din <= x"0208530c";
		wait for Clk_period;
		Addr <=  "0011010110111";
		Trees_din <= x"04022508";
		wait for Clk_period;
		Addr <=  "0011010111000";
		Trees_din <= x"04011c04";
		wait for Clk_period;
		Addr <=  "0011010111001";
		Trees_din <= x"00021bbd";
		wait for Clk_period;
		Addr <=  "0011010111010";
		Trees_din <= x"00d51bbd";
		wait for Clk_period;
		Addr <=  "0011010111011";
		Trees_din <= x"ffcf1bbd";
		wait for Clk_period;
		Addr <=  "0011010111100";
		Trees_din <= x"ff841bbd";
		wait for Clk_period;
		Addr <=  "0011010111101";
		Trees_din <= x"07f75020";
		wait for Clk_period;
		Addr <=  "0011010111110";
		Trees_din <= x"0c00af10";
		wait for Clk_period;
		Addr <=  "0011010111111";
		Trees_din <= x"07f70a08";
		wait for Clk_period;
		Addr <=  "0011011000000";
		Trees_din <= x"000f8604";
		wait for Clk_period;
		Addr <=  "0011011000001";
		Trees_din <= x"ff9b1bbd";
		wait for Clk_period;
		Addr <=  "0011011000010";
		Trees_din <= x"003a1bbd";
		wait for Clk_period;
		Addr <=  "0011011000011";
		Trees_din <= x"1f025b04";
		wait for Clk_period;
		Addr <=  "0011011000100";
		Trees_din <= x"ffdf1bbd";
		wait for Clk_period;
		Addr <=  "0011011000101";
		Trees_din <= x"00af1bbd";
		wait for Clk_period;
		Addr <=  "0011011000110";
		Trees_din <= x"0b007608";
		wait for Clk_period;
		Addr <=  "0011011000111";
		Trees_din <= x"0a004204";
		wait for Clk_period;
		Addr <=  "0011011001000";
		Trees_din <= x"00ef1bbd";
		wait for Clk_period;
		Addr <=  "0011011001001";
		Trees_din <= x"003c1bbd";
		wait for Clk_period;
		Addr <=  "0011011001010";
		Trees_din <= x"0b007e04";
		wait for Clk_period;
		Addr <=  "0011011001011";
		Trees_din <= x"ffa11bbd";
		wait for Clk_period;
		Addr <=  "0011011001100";
		Trees_din <= x"00831bbd";
		wait for Clk_period;
		Addr <=  "0011011001101";
		Trees_din <= x"07f77b0c";
		wait for Clk_period;
		Addr <=  "0011011001110";
		Trees_din <= x"0d000104";
		wait for Clk_period;
		Addr <=  "0011011001111";
		Trees_din <= x"fff81bbd";
		wait for Clk_period;
		Addr <=  "0011011010000";
		Trees_din <= x"14039f04";
		wait for Clk_period;
		Addr <=  "0011011010001";
		Trees_din <= x"ffd91bbd";
		wait for Clk_period;
		Addr <=  "0011011010010";
		Trees_din <= x"ff541bbd";
		wait for Clk_period;
		Addr <=  "0011011010011";
		Trees_din <= x"0b007108";
		wait for Clk_period;
		Addr <=  "0011011010100";
		Trees_din <= x"1f028204";
		wait for Clk_period;
		Addr <=  "0011011010101";
		Trees_din <= x"00191bbd";
		wait for Clk_period;
		Addr <=  "0011011010110";
		Trees_din <= x"ffb51bbd";
		wait for Clk_period;
		Addr <=  "0011011010111";
		Trees_din <= x"06feee04";
		wait for Clk_period;
		Addr <=  "0011011011000";
		Trees_din <= x"000d1bbd";
		wait for Clk_period;
		Addr <=  "0011011011001";
		Trees_din <= x"ffe51bbd";
		wait for Clk_period;
		Addr <=  "0011011011010";
		Trees_din <= x"1e028724";
		wait for Clk_period;
		Addr <=  "0011011011011";
		Trees_din <= x"0900e814";
		wait for Clk_period;
		Addr <=  "0011011011100";
		Trees_din <= x"05f1e00c";
		wait for Clk_period;
		Addr <=  "0011011011101";
		Trees_din <= x"1b027708";
		wait for Clk_period;
		Addr <=  "0011011011110";
		Trees_din <= x"0c00aa04";
		wait for Clk_period;
		Addr <=  "0011011011111";
		Trees_din <= x"00231bbd";
		wait for Clk_period;
		Addr <=  "0011011100000";
		Trees_din <= x"ff821bbd";
		wait for Clk_period;
		Addr <=  "0011011100001";
		Trees_din <= x"00701bbd";
		wait for Clk_period;
		Addr <=  "0011011100010";
		Trees_din <= x"04098204";
		wait for Clk_period;
		Addr <=  "0011011100011";
		Trees_din <= x"00931bbd";
		wait for Clk_period;
		Addr <=  "0011011100100";
		Trees_din <= x"000b1bbd";
		wait for Clk_period;
		Addr <=  "0011011100101";
		Trees_din <= x"1000450c";
		wait for Clk_period;
		Addr <=  "0011011100110";
		Trees_din <= x"0900ed08";
		wait for Clk_period;
		Addr <=  "0011011100111";
		Trees_din <= x"1afb7a04";
		wait for Clk_period;
		Addr <=  "0011011101000";
		Trees_din <= x"ff471bbd";
		wait for Clk_period;
		Addr <=  "0011011101001";
		Trees_din <= x"ffd31bbd";
		wait for Clk_period;
		Addr <=  "0011011101010";
		Trees_din <= x"00201bbd";
		wait for Clk_period;
		Addr <=  "0011011101011";
		Trees_din <= x"006a1bbd";
		wait for Clk_period;
		Addr <=  "0011011101100";
		Trees_din <= x"1401a204";
		wait for Clk_period;
		Addr <=  "0011011101101";
		Trees_din <= x"ff851bbd";
		wait for Clk_period;
		Addr <=  "0011011101110";
		Trees_din <= x"00131bbd";
		wait for Clk_period;
		Addr <=  "0011011101111";
		Trees_din <= x"17039b3c";
		wait for Clk_period;
		Addr <=  "0011011110000";
		Trees_din <= x"1efc9510";
		wait for Clk_period;
		Addr <=  "0011011110001";
		Trees_din <= x"1400fb08";
		wait for Clk_period;
		Addr <=  "0011011110010";
		Trees_din <= x"12008304";
		wait for Clk_period;
		Addr <=  "0011011110011";
		Trees_din <= x"00671c51";
		wait for Clk_period;
		Addr <=  "0011011110100";
		Trees_din <= x"ffbc1c51";
		wait for Clk_period;
		Addr <=  "0011011110101";
		Trees_din <= x"0b009b04";
		wait for Clk_period;
		Addr <=  "0011011110110";
		Trees_din <= x"ff5e1c51";
		wait for Clk_period;
		Addr <=  "0011011110111";
		Trees_din <= x"ffd01c51";
		wait for Clk_period;
		Addr <=  "0011011111000";
		Trees_din <= x"08005020";
		wait for Clk_period;
		Addr <=  "0011011111001";
		Trees_din <= x"21002510";
		wait for Clk_period;
		Addr <=  "0011011111010";
		Trees_din <= x"20040008";
		wait for Clk_period;
		Addr <=  "0011011111011";
		Trees_din <= x"07f83c04";
		wait for Clk_period;
		Addr <=  "0011011111100";
		Trees_din <= x"00811c51";
		wait for Clk_period;
		Addr <=  "0011011111101";
		Trees_din <= x"ff881c51";
		wait for Clk_period;
		Addr <=  "0011011111110";
		Trees_din <= x"21000004";
		wait for Clk_period;
		Addr <=  "0011011111111";
		Trees_din <= x"00001c51";
		wait for Clk_period;
		Addr <=  "0011100000000";
		Trees_din <= x"00391c51";
		wait for Clk_period;
		Addr <=  "0011100000001";
		Trees_din <= x"010d1608";
		wait for Clk_period;
		Addr <=  "0011100000010";
		Trees_din <= x"0b007704";
		wait for Clk_period;
		Addr <=  "0011100000011";
		Trees_din <= x"ffdd1c51";
		wait for Clk_period;
		Addr <=  "0011100000100";
		Trees_din <= x"00791c51";
		wait for Clk_period;
		Addr <=  "0011100000101";
		Trees_din <= x"12008904";
		wait for Clk_period;
		Addr <=  "0011100000110";
		Trees_din <= x"ff911c51";
		wait for Clk_period;
		Addr <=  "0011100000111";
		Trees_din <= x"002e1c51";
		wait for Clk_period;
		Addr <=  "0011100001000";
		Trees_din <= x"21000008";
		wait for Clk_period;
		Addr <=  "0011100001001";
		Trees_din <= x"0c00c504";
		wait for Clk_period;
		Addr <=  "0011100001010";
		Trees_din <= x"00231c51";
		wait for Clk_period;
		Addr <=  "0011100001011";
		Trees_din <= x"00e41c51";
		wait for Clk_period;
		Addr <=  "0011100001100";
		Trees_din <= x"ff981c51";
		wait for Clk_period;
		Addr <=  "0011100001101";
		Trees_din <= x"000a8804";
		wait for Clk_period;
		Addr <=  "0011100001110";
		Trees_din <= x"ffde1c51";
		wait for Clk_period;
		Addr <=  "0011100001111";
		Trees_din <= x"0c00c108";
		wait for Clk_period;
		Addr <=  "0011100010000";
		Trees_din <= x"02073804";
		wait for Clk_period;
		Addr <=  "0011100010001";
		Trees_din <= x"00e61c51";
		wait for Clk_period;
		Addr <=  "0011100010010";
		Trees_din <= x"002a1c51";
		wait for Clk_period;
		Addr <=  "0011100010011";
		Trees_din <= x"ffff1c51";
		wait for Clk_period;
		Addr <=  "0011100010100";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  2
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"07072364";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"0703c338";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"0701e41c";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"07ff5c0c";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"11038704";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"ff520125";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"09006704";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"00370125";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"ff770125";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"1400e308";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"00053f04";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"ff840125";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"00ca0125";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"08004c04";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"ff610125";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"ffc70125";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"0600050c";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"22000108";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"02051304";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"ff550125";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"ff950125";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"000f0125";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"03f9d108";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"12006e04";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"005f0125";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"ff600125";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"08004204";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"ff9c0125";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"01ca0125";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"010dbd1c";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"0b008c10";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"04facb08";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"0e003f04";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"ff630125";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"00df0125";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"10004604";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"001f0125";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"01870125";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"01008904";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"ffa40125";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"1afc4804";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"02c70125";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"00890125";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"1101a904";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"ff5a0125";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"16006108";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"03f90904";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"ff960125";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"015c0125";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"ff650125";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"010c9118";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"0301e210";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"0006db0c";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"010a6404";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"03ff0125";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"010ac004";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"00890125";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"02a80125";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"00df0125";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"00fef404";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"00370125";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"015c0125";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"070b480c";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"00049608";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"17f71104";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"00000125";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"ff620125";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"00c20125";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"0e002c04";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"ffa40125";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"0d005804";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"00ca0125";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"02e70125";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"0706185c";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"0703c338";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"0701e41c";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"07ff5c0c";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"13008808";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"01050e04";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"003a0249";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"ff820249";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"ff580249";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"1400e308";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"0900bc04";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"ff8a0249";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"00d80249";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"0900ef04";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"ff650249";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"ffb10249";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"0600050c";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"22000108";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"19000b04";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"ff620249";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"ffbc0249";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"00160249";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"10004c08";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"04fe2a04";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"ff660249";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"00140249";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"0b007604";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"01440249";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"ff8f0249";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"06fdee10";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"11000204";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"00d20249";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"0c00b204";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"ff5f0249";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"0900da04";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"ff8c0249";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"009a0249";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"03fc1e10";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"1c025b08";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"04fc7e04";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"ff8b0249";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"01ce0249";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"0a004204";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"00340249";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"ff820249";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"01e10249";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"010c9120";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"03f55108";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"0d00e004";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"ff950249";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"00c50249";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"1300f408";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"00ff1204";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"ff930249";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"01160249";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"19001708";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"10004704";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"015c0249";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"01e00249";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"15003a04";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"01510249";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"ff7a0249";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"070b4810";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"03f62904";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"00da0249";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"08004504";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"ff630249";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"0200b504";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"00b40249";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"ff840249";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"0e002c04";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"ffa60249";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"01930249";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"0705714c";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"0701e424";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"07ff5c0c";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"11038704";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"ff5c0355";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"0c00aa04";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"ff8b0355";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"003f0355";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"1400e308";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"010d9f04";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"ff8e0355";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"00d00355";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"0900ef08";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"08004c04";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"ff650355";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"ffef0355";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"12007504";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"ff800355";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"00eb0355";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"010dbd1c";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"0e004510";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"0703c308";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"0a004604";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"ff7c0355";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"fff20355";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"19000604";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"ffeb0355";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"00c50355";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"05f57d04";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"ffa70355";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"06fe0e04";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"001e0355";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"01930355";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"05f20e08";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"0a004004";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"00420355";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"ff970355";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"ff5f0355";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"010b2818";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"050b6014";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"0307c210";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"06ff3108";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"19001704";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"013c0355";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"00880355";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"10004304";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"00030355";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"012b0355";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"ffa30355";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"ffa20355";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"070b4814";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"04fa5508";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"0e001b04";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"00300355";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"ff610355";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"15003704";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"ff740355";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"0111b004";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"00ee0355";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"ff940355";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"01105f0c";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"03ff7308";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"05f78604";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"018d0355";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"00240355";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"001d0355";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"00040355";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"07057148";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"0701e424";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"07ff5c0c";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"13008808";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"05f7eb04";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"ff930471";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"00400471";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"ff5f0471";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"1400e308";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"00053f04";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"ff950471";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"00b80471";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"0f000808";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"16005904";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"009b0471";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"ff8e0471";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"2003ff04";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"fffa0471";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"ff5e0471";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"010dbd18";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"0e004510";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"06fe0908";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"0704e004";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"ff800471";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"007b0471";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"06fe6604";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"011c0471";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"ffea0471";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"05f67504";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"fff30471";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"010b0471";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"05f20e08";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"12007a04";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"ffa00471";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"00410471";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"ff630471";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"010f713c";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"070a0720";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"05f5f610";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"0d02d108";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"0b008004";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"ff520471";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"00510471";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"05f40e04";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"014e0471";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"00190471";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"03f6b008";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"12007104";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"00240471";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"ff6b0471";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"04fa0c04";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"00140471";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"00e70471";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"04fad710";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"070c0a08";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"03f83904";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"ff610471";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"007f0471";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"0a005004";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"010b0471";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"003d0471";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"1102cb08";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"06f8fa04";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"00510471";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"012a0471";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"00730471";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"15004d08";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"0705b804";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"00670471";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"ff690471";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"00d10471";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"0703c32c";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"07ff5c0c";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"11038704";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"ff61056d";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"10005304";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"ff9f056d";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"0042056d";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"2100681c";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"0600100c";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"07ff6f04";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"002b056d";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"0b00bd04";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"ff76056d";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"0033056d";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"0600ea08";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"08004104";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"ffa2056d";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"00b9056d";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"11031404";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"ff80056d";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"0085056d";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"0091056d";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"07086d30";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"010e111c";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"0c00ce10";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"0f000608";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"03f6e904";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"ffb3056d";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"00c2056d";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"05fb9604";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"ffb9056d";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"0070056d";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"04f9f604";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"ffeb056d";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"15003004";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"0076056d";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"0149056d";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"1101a904";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"ff6c056d";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"0900e008";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"14036904";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"002a056d";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"ff7f056d";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"1403d604";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"003a056d";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"00db056d";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"01105f1c";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"070c0a10";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"06f95808";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"0e004404";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"ff5e056d";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"0086056d";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"06005d04";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"00b6056d";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"002c056d";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"04fd3808";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"1600a304";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"00e9056d";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"0033056d";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"0045056d";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"1afbca04";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"002f056d";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"ff9c056d";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"0703c330";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"07ff5c0c";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"11038704";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"ff640691";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"0205a804";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"00400691";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"ffa50691";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"21006820";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"06001010";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"0e002808";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"15003904";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"ff930691";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"005d0691";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"00fcb404";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"ffe10691";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"ff690691";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"06009308";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"1afcc004";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"00940691";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"ff950691";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"07024804";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"ff7e0691";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"001c0691";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"00820691";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"070a0738";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"05f56318";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"12008810";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"0d02eb08";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"00200691";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"ff550691";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"10004a04";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"00e00691";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"ff990691";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"0204bf04";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"ffa10691";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"00fa0691";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"04fa0c10";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"0d000008";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"0a004504";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"00e80691";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"00460691";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"00fbbc04";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"00810691";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"ff990691";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"0900e808";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"03f6b004";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"ffc20691";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"00bf0691";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"0a003d04";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"00be0691";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"ff8c0691";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"04fad71c";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"070c0a0c";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"12006f04";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"00c80691";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"10004404";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"005a0691";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"ff6f0691";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"0a005008";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"03f9ea04";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"00690691";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"00d60691";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"02fed204";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"008f0691";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"ff810691";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"04fe3708";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"0f013e04";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"00e80691";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"00290691";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"19000004";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"ffb30691";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"00b40691";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"0703c338";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"07ff5c18";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"13008804";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"fff507c5";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"12005a08";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"1303bb04";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"004807c5";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"ff7d07c5";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"04f9de08";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"0c00cd04";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"ff7b07c5";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"004807c5";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"ff6307c5";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"2100681c";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"0900ef10";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"0900c308";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"0900bc04";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"ffa707c5";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"008c07c5";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"0a003b04";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"000007c5";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"ff6207c5";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"0c00a608";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"0206d504";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"ff7207c5";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"007a07c5";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"012907c5";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"007407c5";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"070a0738";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"05f56318";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"12008810";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"0d02eb08";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"002307c5";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"ff5907c5";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"10004a04";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"00d007c5";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"ff9f07c5";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"0204bf04";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"ffa907c5";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"00d407c5";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"04fa0c10";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"1303a908";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"10005304";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"ff5b07c5";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"001307c5";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"05f90204";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"ffba07c5";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"00b607c5";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"03f6b008";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"0d025604";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"ff6407c5";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"00b207c5";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"0900e804";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"009f07c5";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"fff407c5";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"04fad71c";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"070c0a0c";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"12006f04";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"00b107c5";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"10004404";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"004b07c5";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"ff7907c5";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"0a005008";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"18001d04";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"005707c5";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"00c207c5";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"02fed204";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"008307c5";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"ff8407c5";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"1102cb0c";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"0600e108";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"06f8fa04";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"002907c5";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"00d707c5";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"002107c5";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"002e07c5";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"0703c334";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"07ff5c18";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"11038714";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"12005a08";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"0e004304";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"004908cd";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"ff8108cd";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"04f9de08";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"15003204";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"004808cd";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"ff8108cd";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"ff6508cd";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"fffe08cd";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"02021704";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"ff6a08cd";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"05fc130c";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"2003fb04";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"008008cd";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"1400e304";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"005c08cd";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"ffa508cd";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"18001604";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"014e08cd";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"09009804";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"006908cd";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"ff7b08cd";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"070c0a38";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"03f8ba20";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"1403f610";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"04fc1d08";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"0a003c04";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"007808cd";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"ff8008cd";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"1101b304";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"001208cd";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"00ea08cd";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"17f74208";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"01077704";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"009008cd";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"ff8f08cd";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"0a003c04";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"005c08cd";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"ff5708cd";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"02064e10";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"0900e708";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"1303d904";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"003e08cd";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"00c208cd";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"00ff1204";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"008208cd";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"ffb008cd";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"0705de04";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"ff7608cd";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"000908cd";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"08004414";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"010a640c";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"1afae208";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"1c028404";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"ff9b08cd";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"008f08cd";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"00b208cd";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"010f1504";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"ff7208cd";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"004808cd";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"00c508cd";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"07024844";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"07fef110";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"13008804";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"000c0a11";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"12005a08";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"0e004304";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"004a0a11";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"ff860a11";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"ff660a11";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"12007b18";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"0e00410c";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"14040004";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"ff660a11";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"0900f104";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"ff8f0a11";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"00450a11";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"08004508";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"12005f04";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"ff970a11";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"00db0a11";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"ff7e0a11";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"0007370c";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"17f79808";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"06fefa04";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"ff900a11";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"00ae0a11";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"ff6c0a11";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"10004108";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"06ff2004";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"ff8c0a11";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"00440a11";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"0b008404";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"014c0a11";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"00070a11";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"070a0738";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"05f56818";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"0b00860c";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"05f39208";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"03fa4604";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"ff720a11";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"00800a11";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"ff610a11";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"010e1108";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"10003d04";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"000d0a11";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"00e30a11";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"ff9a0a11";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"19000810";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"12007408";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"010b8304";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"008a0a11";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"ffbb0a11";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"07040e04";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"ff6d0a11";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"000c0a11";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"1e028508";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"17f8bd04";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"007e0a11";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"ffb30a11";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"1afea704";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"01430a11";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"00670a11";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"04fad718";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"070c0a0c";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"12006f04";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"00920a11";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"12007504";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"ff670a11";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"00250a11";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"08004408";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"010a6404";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"00840a11";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"ffab0a11";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"00b60a11";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"04fe3708";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"0f013e04";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"00bf0a11";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"000d0a11";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"08003f04";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"ffa70a11";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"00830a11";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"0702483c";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"07fef118";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"11038714";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"12005a08";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"11008804";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"ff8b0b4d";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"00490b4d";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"1d028604";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"ff650b4d";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"0209ab04";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"ff7c0b4d";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"00450b4d";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"00110b4d";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"0a003d0c";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"08004004";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"ff880b4d";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"1100fb04";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"01de0b4d";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"ffa60b4d";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"08004c10";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"0900ef08";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"0d02bf04";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"ff810b4d";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"00070b4d";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"12007504";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"ff850b4d";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"00d40b4d";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"18007904";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"00db0b4d";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"ffa20b4d";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"070a0734";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"05f56818";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"0b00860c";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"05f39208";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"0d011b04";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"ff780b4d";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"007f0b4d";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"ff650b4d";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"010b8304";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"00b30b4d";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"11016a04";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"ff9d0b4d";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"00230b4d";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"19000810";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"12007408";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"010c5204";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"006f0b4d";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"ffb10b4d";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"19000204";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"00090b4d";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"ff600b4d";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"04fa3304";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"ffb60b4d";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"05039704";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"00d90b4d";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"ffaa0b4d";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"04fab720";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"1c027510";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"010a9f08";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"0900ef04";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"00a20b4d";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"fff60b4d";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"0900bc04";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"ffc30b4d";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"007f0b4d";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"04f8d408";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"0b006d04";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"fff40b4d";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"00850b4d";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"08004604";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"ff4f0b4d";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"00180b4d";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"1102cb08";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"06f8fa04";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"00160b4d";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"00b00b4d";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"06fd6e04";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"00600b4d";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"ff9f0b4d";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"0701e43c";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"07fe6614";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"03fc760c";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"1d028604";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"ff660c31";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"0209ab04";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"ff820c31";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"00430c31";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"05f61a04";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"004b0c31";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"ff930c31";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"1100fb1c";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"1e02620c";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"0e004104";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"ff700c31";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"0e004404";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"00c40c31";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"ff980c31";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"1b026708";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"16006a04";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"01320c31";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"ffb10c31";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"1100da04";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"ff7b0c31";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"009e0c31";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"04008e04";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"ff6a0c31";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"02043b04";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"00c60c31";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"ff9f0c31";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"070c0a20";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"02fe920c";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"0d001504";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"00250c31";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"1b025a04";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"ffd10c31";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"ff4d0c31";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"0111b010";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"0900e008";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"05f33104";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"ff7d0c31";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"00440c31";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"16006004";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"ff860c31";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"001a0c31";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"ff860c31";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"08004414";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"010a640c";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"1afae208";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"1c028404";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"ff9e0c31";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"00720c31";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"00980c31";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"04f9de04";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"ff850c31";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"00440c31";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"00a90c31";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"0701e43c";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"07fe6614";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"12005a08";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"0205a804";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"00490d4d";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"ff9a0d4d";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"0606cc04";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"ff660d4d";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"11024004";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"ff860d4d";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"00480d4d";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"0a003d0c";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"08004004";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"ff930d4d";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"1303a004";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"fff60d4d";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"016a0d4d";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"0b007d0c";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"11002108";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"0000f704";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"00b40d4d";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"ff890d4d";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"ff6a0d4d";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"0b008408";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"10004104";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"ffa60d4d";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"00bb0d4d";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"10005304";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"ff730d4d";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"00580d4d";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"07061834";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"06fdee14";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"0900db08";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"0200d204";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"fff10d4d";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"ff630d4d";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"06fc5f08";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"0e002b04";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"00990d4d";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"ffce0d4d";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"ff8c0d4d";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"15003b10";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"06fe3e08";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"1e027404";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"002a0d4d";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"00d00d4d";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"1e028704";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"ff8a0d4d";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"00590d4d";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"0e003808";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"03f66c04";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"ffde0d4d";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"00b90d4d";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"03fa9504";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"ffa70d4d";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"008c0d4d";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"01023408";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"03f62904";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"00060d4d";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"00a70d4d";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"06ff310c";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"1300b204";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"ff820d4d";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"1b024604";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"ffe00d4d";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"00570d4d";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"0a003d04";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"00800d4d";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"0201b104";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"ff640d4d";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"fffd0d4d";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"07002028";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"0a005a20";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"04fc120c";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"0b005e04";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"00860e51";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"0f010c04";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"ff770e51";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"00420e51";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"06fb8b08";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"15003a04";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"004a0e51";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"ffad0e51";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"1d028604";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"ff670e51";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"14039f04";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"ff8a0e51";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"00460e51";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"03fa5f04";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"ffa00e51";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"009d0e51";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"0703c330";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"0900ef20";
		wait for Clk_period;
		Addr <=  "0001101101001";
		Trees_din <= x"09009910";
		wait for Clk_period;
		Addr <=  "0001101101010";
		Trees_din <= x"0a004e08";
		wait for Clk_period;
		Addr <=  "0001101101011";
		Trees_din <= x"05f6d304";
		wait for Clk_period;
		Addr <=  "0001101101100";
		Trees_din <= x"ff9a0e51";
		wait for Clk_period;
		Addr <=  "0001101101101";
		Trees_din <= x"00c20e51";
		wait for Clk_period;
		Addr <=  "0001101101110";
		Trees_din <= x"0e003d04";
		wait for Clk_period;
		Addr <=  "0001101101111";
		Trees_din <= x"ff7b0e51";
		wait for Clk_period;
		Addr <=  "0001101110000";
		Trees_din <= x"005e0e51";
		wait for Clk_period;
		Addr <=  "0001101110001";
		Trees_din <= x"12006e08";
		wait for Clk_period;
		Addr <=  "0001101110010";
		Trees_din <= x"00050704";
		wait for Clk_period;
		Addr <=  "0001101110011";
		Trees_din <= x"00500e51";
		wait for Clk_period;
		Addr <=  "0001101110100";
		Trees_din <= x"ff900e51";
		wait for Clk_period;
		Addr <=  "0001101110101";
		Trees_din <= x"07004504";
		wait for Clk_period;
		Addr <=  "0001101110110";
		Trees_din <= x"00420e51";
		wait for Clk_period;
		Addr <=  "0001101110111";
		Trees_din <= x"ff770e51";
		wait for Clk_period;
		Addr <=  "0001101111000";
		Trees_din <= x"0c009808";
		wait for Clk_period;
		Addr <=  "0001101111001";
		Trees_din <= x"1f024804";
		wait for Clk_period;
		Addr <=  "0001101111010";
		Trees_din <= x"00340e51";
		wait for Clk_period;
		Addr <=  "0001101111011";
		Trees_din <= x"ff8e0e51";
		wait for Clk_period;
		Addr <=  "0001101111100";
		Trees_din <= x"02062604";
		wait for Clk_period;
		Addr <=  "0001101111101";
		Trees_din <= x"00020e51";
		wait for Clk_period;
		Addr <=  "0001101111110";
		Trees_din <= x"011d0e51";
		wait for Clk_period;
		Addr <=  "0001101111111";
		Trees_din <= x"070c0a1c";
		wait for Clk_period;
		Addr <=  "0001110000000";
		Trees_din <= x"0c00d610";
		wait for Clk_period;
		Addr <=  "0001110000001";
		Trees_din <= x"04faec08";
		wait for Clk_period;
		Addr <=  "0001110000010";
		Trees_din <= x"0d006504";
		wait for Clk_period;
		Addr <=  "0001110000011";
		Trees_din <= x"00210e51";
		wait for Clk_period;
		Addr <=  "0001110000100";
		Trees_din <= x"ff8e0e51";
		wait for Clk_period;
		Addr <=  "0001110000101";
		Trees_din <= x"02031b04";
		wait for Clk_period;
		Addr <=  "0001110000110";
		Trees_din <= x"00610e51";
		wait for Clk_period;
		Addr <=  "0001110000111";
		Trees_din <= x"fff00e51";
		wait for Clk_period;
		Addr <=  "0001110001000";
		Trees_din <= x"06fb6204";
		wait for Clk_period;
		Addr <=  "0001110001001";
		Trees_din <= x"ffbd0e51";
		wait for Clk_period;
		Addr <=  "0001110001010";
		Trees_din <= x"1403fe04";
		wait for Clk_period;
		Addr <=  "0001110001011";
		Trees_din <= x"00a20e51";
		wait for Clk_period;
		Addr <=  "0001110001100";
		Trees_din <= x"ffd90e51";
		wait for Clk_period;
		Addr <=  "0001110001101";
		Trees_din <= x"0800440c";
		wait for Clk_period;
		Addr <=  "0001110001110";
		Trees_din <= x"0900e108";
		wait for Clk_period;
		Addr <=  "0001110001111";
		Trees_din <= x"05f77a04";
		wait for Clk_period;
		Addr <=  "0001110010000";
		Trees_din <= x"ffb10e51";
		wait for Clk_period;
		Addr <=  "0001110010001";
		Trees_din <= x"004b0e51";
		wait for Clk_period;
		Addr <=  "0001110010010";
		Trees_din <= x"00890e51";
		wait for Clk_period;
		Addr <=  "0001110010011";
		Trees_din <= x"009c0e51";
		wait for Clk_period;
		Addr <=  "0001110010100";
		Trees_din <= x"07fef114";
		wait for Clk_period;
		Addr <=  "0001110010101";
		Trees_din <= x"0005d210";
		wait for Clk_period;
		Addr <=  "0001110010110";
		Trees_din <= x"0003e304";
		wait for Clk_period;
		Addr <=  "0001110010111";
		Trees_din <= x"ff7a0f25";
		wait for Clk_period;
		Addr <=  "0001110011000";
		Trees_din <= x"18008a04";
		wait for Clk_period;
		Addr <=  "0001110011001";
		Trees_din <= x"ff9a0f25";
		wait for Clk_period;
		Addr <=  "0001110011010";
		Trees_din <= x"08003f04";
		wait for Clk_period;
		Addr <=  "0001110011011";
		Trees_din <= x"010b0f25";
		wait for Clk_period;
		Addr <=  "0001110011100";
		Trees_din <= x"ffae0f25";
		wait for Clk_period;
		Addr <=  "0001110011101";
		Trees_din <= x"ff680f25";
		wait for Clk_period;
		Addr <=  "0001110011110";
		Trees_din <= x"0703c324";
		wait for Clk_period;
		Addr <=  "0001110011111";
		Trees_din <= x"02021704";
		wait for Clk_period;
		Addr <=  "0001110100000";
		Trees_din <= x"ff740f25";
		wait for Clk_period;
		Addr <=  "0001110100001";
		Trees_din <= x"0109bb10";
		wait for Clk_period;
		Addr <=  "0001110100010";
		Trees_din <= x"1403ff08";
		wait for Clk_period;
		Addr <=  "0001110100011";
		Trees_din <= x"0900f004";
		wait for Clk_period;
		Addr <=  "0001110100100";
		Trees_din <= x"ff7d0f25";
		wait for Clk_period;
		Addr <=  "0001110100101";
		Trees_din <= x"00300f25";
		wait for Clk_period;
		Addr <=  "0001110100110";
		Trees_din <= x"0f000204";
		wait for Clk_period;
		Addr <=  "0001110100111";
		Trees_din <= x"ff960f25";
		wait for Clk_period;
		Addr <=  "0001110101000";
		Trees_din <= x"00700f25";
		wait for Clk_period;
		Addr <=  "0001110101001";
		Trees_din <= x"12008108";
		wait for Clk_period;
		Addr <=  "0001110101010";
		Trees_din <= x"010b8304";
		wait for Clk_period;
		Addr <=  "0001110101011";
		Trees_din <= x"00410f25";
		wait for Clk_period;
		Addr <=  "0001110101100";
		Trees_din <= x"ff900f25";
		wait for Clk_period;
		Addr <=  "0001110101101";
		Trees_din <= x"0b008304";
		wait for Clk_period;
		Addr <=  "0001110101110";
		Trees_din <= x"01610f25";
		wait for Clk_period;
		Addr <=  "0001110101111";
		Trees_din <= x"00040f25";
		wait for Clk_period;
		Addr <=  "0001110110000";
		Trees_din <= x"03f8f520";
		wait for Clk_period;
		Addr <=  "0001110110001";
		Trees_din <= x"0d00aa10";
		wait for Clk_period;
		Addr <=  "0001110110010";
		Trees_din <= x"1c026208";
		wait for Clk_period;
		Addr <=  "0001110110011";
		Trees_din <= x"0705b804";
		wait for Clk_period;
		Addr <=  "0001110110100";
		Trees_din <= x"ff970f25";
		wait for Clk_period;
		Addr <=  "0001110110101";
		Trees_din <= x"005e0f25";
		wait for Clk_period;
		Addr <=  "0001110110110";
		Trees_din <= x"22000004";
		wait for Clk_period;
		Addr <=  "0001110110111";
		Trees_din <= x"ff590f25";
		wait for Clk_period;
		Addr <=  "0001110111000";
		Trees_din <= x"ffef0f25";
		wait for Clk_period;
		Addr <=  "0001110111001";
		Trees_din <= x"04fd3008";
		wait for Clk_period;
		Addr <=  "0001110111010";
		Trees_din <= x"0f003304";
		wait for Clk_period;
		Addr <=  "0001110111011";
		Trees_din <= x"ffae0f25";
		wait for Clk_period;
		Addr <=  "0001110111100";
		Trees_din <= x"00790f25";
		wait for Clk_period;
		Addr <=  "0001110111101";
		Trees_din <= x"11012f04";
		wait for Clk_period;
		Addr <=  "0001110111110";
		Trees_din <= x"fff80f25";
		wait for Clk_period;
		Addr <=  "0001110111111";
		Trees_din <= x"00a90f25";
		wait for Clk_period;
		Addr <=  "0001111000000";
		Trees_din <= x"02064e10";
		wait for Clk_period;
		Addr <=  "0001111000001";
		Trees_din <= x"0d015b08";
		wait for Clk_period;
		Addr <=  "0001111000010";
		Trees_din <= x"0900e704";
		wait for Clk_period;
		Addr <=  "0001111000011";
		Trees_din <= x"00790f25";
		wait for Clk_period;
		Addr <=  "0001111000100";
		Trees_din <= x"fffd0f25";
		wait for Clk_period;
		Addr <=  "0001111000101";
		Trees_din <= x"0d030104";
		wait for Clk_period;
		Addr <=  "0001111000110";
		Trees_din <= x"ffc30f25";
		wait for Clk_period;
		Addr <=  "0001111000111";
		Trees_din <= x"00640f25";
		wait for Clk_period;
		Addr <=  "0001111001000";
		Trees_din <= x"ff730f25";
		wait for Clk_period;
		Addr <=  "0001111001001";
		Trees_din <= x"07fef114";
		wait for Clk_period;
		Addr <=  "0001111001010";
		Trees_din <= x"0005d210";
		wait for Clk_period;
		Addr <=  "0001111001011";
		Trees_din <= x"05f61a08";
		wait for Clk_period;
		Addr <=  "0001111001100";
		Trees_din <= x"0900db04";
		wait for Clk_period;
		Addr <=  "0001111001101";
		Trees_din <= x"ffa80fe9";
		wait for Clk_period;
		Addr <=  "0001111001110";
		Trees_din <= x"00d40fe9";
		wait for Clk_period;
		Addr <=  "0001111001111";
		Trees_din <= x"09006704";
		wait for Clk_period;
		Addr <=  "0001111010000";
		Trees_din <= x"001e0fe9";
		wait for Clk_period;
		Addr <=  "0001111010001";
		Trees_din <= x"ff7b0fe9";
		wait for Clk_period;
		Addr <=  "0001111010010";
		Trees_din <= x"ff690fe9";
		wait for Clk_period;
		Addr <=  "0001111010011";
		Trees_din <= x"0703c324";
		wait for Clk_period;
		Addr <=  "0001111010100";
		Trees_din <= x"02021704";
		wait for Clk_period;
		Addr <=  "0001111010101";
		Trees_din <= x"ff780fe9";
		wait for Clk_period;
		Addr <=  "0001111010110";
		Trees_din <= x"0109bb10";
		wait for Clk_period;
		Addr <=  "0001111010111";
		Trees_din <= x"0f000808";
		wait for Clk_period;
		Addr <=  "0001111011000";
		Trees_din <= x"05f6e204";
		wait for Clk_period;
		Addr <=  "0001111011001";
		Trees_din <= x"ff8e0fe9";
		wait for Clk_period;
		Addr <=  "0001111011010";
		Trees_din <= x"00660fe9";
		wait for Clk_period;
		Addr <=  "0001111011011";
		Trees_din <= x"0900f004";
		wait for Clk_period;
		Addr <=  "0001111011100";
		Trees_din <= x"ff7a0fe9";
		wait for Clk_period;
		Addr <=  "0001111011101";
		Trees_din <= x"00210fe9";
		wait for Clk_period;
		Addr <=  "0001111011110";
		Trees_din <= x"12008108";
		wait for Clk_period;
		Addr <=  "0001111011111";
		Trees_din <= x"010b8304";
		wait for Clk_period;
		Addr <=  "0001111100000";
		Trees_din <= x"00360fe9";
		wait for Clk_period;
		Addr <=  "0001111100001";
		Trees_din <= x"ff960fe9";
		wait for Clk_period;
		Addr <=  "0001111100010";
		Trees_din <= x"0b008304";
		wait for Clk_period;
		Addr <=  "0001111100011";
		Trees_din <= x"010e0fe9";
		wait for Clk_period;
		Addr <=  "0001111100100";
		Trees_din <= x"00070fe9";
		wait for Clk_period;
		Addr <=  "0001111100101";
		Trees_din <= x"070c0a18";
		wait for Clk_period;
		Addr <=  "0001111100110";
		Trees_din <= x"02fe9208";
		wait for Clk_period;
		Addr <=  "0001111100111";
		Trees_din <= x"17f82e04";
		wait for Clk_period;
		Addr <=  "0001111101000";
		Trees_din <= x"ff6a0fe9";
		wait for Clk_period;
		Addr <=  "0001111101001";
		Trees_din <= x"001c0fe9";
		wait for Clk_period;
		Addr <=  "0001111101010";
		Trees_din <= x"0900e708";
		wait for Clk_period;
		Addr <=  "0001111101011";
		Trees_din <= x"17f72204";
		wait for Clk_period;
		Addr <=  "0001111101100";
		Trees_din <= x"00a10fe9";
		wait for Clk_period;
		Addr <=  "0001111101101";
		Trees_din <= x"001a0fe9";
		wait for Clk_period;
		Addr <=  "0001111101110";
		Trees_din <= x"01077704";
		wait for Clk_period;
		Addr <=  "0001111101111";
		Trees_din <= x"00430fe9";
		wait for Clk_period;
		Addr <=  "0001111110000";
		Trees_din <= x"ff8f0fe9";
		wait for Clk_period;
		Addr <=  "0001111110001";
		Trees_din <= x"0f00370c";
		wait for Clk_period;
		Addr <=  "0001111110010";
		Trees_din <= x"1403ff04";
		wait for Clk_period;
		Addr <=  "0001111110011";
		Trees_din <= x"008d0fe9";
		wait for Clk_period;
		Addr <=  "0001111110100";
		Trees_din <= x"17f77a04";
		wait for Clk_period;
		Addr <=  "0001111110101";
		Trees_din <= x"00730fe9";
		wait for Clk_period;
		Addr <=  "0001111110110";
		Trees_din <= x"ffa70fe9";
		wait for Clk_period;
		Addr <=  "0001111110111";
		Trees_din <= x"0b007c04";
		wait for Clk_period;
		Addr <=  "0001111111000";
		Trees_din <= x"005a0fe9";
		wait for Clk_period;
		Addr <=  "0001111111001";
		Trees_din <= x"ffb70fe9";
		wait for Clk_period;
		Addr <=  "0001111111010";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0001111111011";
		Trees_din <= x"07fef114";
		wait for Clk_period;
		Addr <=  "0001111111100";
		Trees_din <= x"0005d210";
		wait for Clk_period;
		Addr <=  "0001111111101";
		Trees_din <= x"0003e304";
		wait for Clk_period;
		Addr <=  "0001111111110";
		Trees_din <= x"ff8110a1";
		wait for Clk_period;
		Addr <=  "0001111111111";
		Trees_din <= x"1303bb08";
		wait for Clk_period;
		Addr <=  "0010000000000";
		Trees_din <= x"05f65604";
		wait for Clk_period;
		Addr <=  "0010000000001";
		Trees_din <= x"00e310a1";
		wait for Clk_period;
		Addr <=  "0010000000010";
		Trees_din <= x"fffb10a1";
		wait for Clk_period;
		Addr <=  "0010000000011";
		Trees_din <= x"ff9f10a1";
		wait for Clk_period;
		Addr <=  "0010000000100";
		Trees_din <= x"ff6a10a1";
		wait for Clk_period;
		Addr <=  "0010000000101";
		Trees_din <= x"070c0a34";
		wait for Clk_period;
		Addr <=  "0010000000110";
		Trees_din <= x"0c00dc18";
		wait for Clk_period;
		Addr <=  "0010000000111";
		Trees_din <= x"22000510";
		wait for Clk_period;
		Addr <=  "0010000001000";
		Trees_din <= x"04faec08";
		wait for Clk_period;
		Addr <=  "0010000001001";
		Trees_din <= x"0d006504";
		wait for Clk_period;
		Addr <=  "0010000001010";
		Trees_din <= x"fff810a1";
		wait for Clk_period;
		Addr <=  "0010000001011";
		Trees_din <= x"ff8f10a1";
		wait for Clk_period;
		Addr <=  "0010000001100";
		Trees_din <= x"03fa3904";
		wait for Clk_period;
		Addr <=  "0010000001101";
		Trees_din <= x"ffe810a1";
		wait for Clk_period;
		Addr <=  "0010000001110";
		Trees_din <= x"003b10a1";
		wait for Clk_period;
		Addr <=  "0010000001111";
		Trees_din <= x"22000a04";
		wait for Clk_period;
		Addr <=  "0010000010000";
		Trees_din <= x"00c910a1";
		wait for Clk_period;
		Addr <=  "0010000010001";
		Trees_din <= x"001710a1";
		wait for Clk_period;
		Addr <=  "0010000010010";
		Trees_din <= x"12009710";
		wait for Clk_period;
		Addr <=  "0010000010011";
		Trees_din <= x"18006608";
		wait for Clk_period;
		Addr <=  "0010000010100";
		Trees_din <= x"0e001e04";
		wait for Clk_period;
		Addr <=  "0010000010101";
		Trees_din <= x"002810a1";
		wait for Clk_period;
		Addr <=  "0010000010110";
		Trees_din <= x"ffaa10a1";
		wait for Clk_period;
		Addr <=  "0010000010111";
		Trees_din <= x"19000d04";
		wait for Clk_period;
		Addr <=  "0010000011000";
		Trees_din <= x"00d410a1";
		wait for Clk_period;
		Addr <=  "0010000011001";
		Trees_din <= x"002610a1";
		wait for Clk_period;
		Addr <=  "0010000011010";
		Trees_din <= x"0002ed08";
		wait for Clk_period;
		Addr <=  "0010000011011";
		Trees_din <= x"03f84a04";
		wait for Clk_period;
		Addr <=  "0010000011100";
		Trees_din <= x"005d10a1";
		wait for Clk_period;
		Addr <=  "0010000011101";
		Trees_din <= x"fff510a1";
		wait for Clk_period;
		Addr <=  "0010000011110";
		Trees_din <= x"ff8810a1";
		wait for Clk_period;
		Addr <=  "0010000011111";
		Trees_din <= x"08003a08";
		wait for Clk_period;
		Addr <=  "0010000100000";
		Trees_din <= x"1c025104";
		wait for Clk_period;
		Addr <=  "0010000100001";
		Trees_din <= x"006410a1";
		wait for Clk_period;
		Addr <=  "0010000100010";
		Trees_din <= x"ffa710a1";
		wait for Clk_period;
		Addr <=  "0010000100011";
		Trees_din <= x"1303d404";
		wait for Clk_period;
		Addr <=  "0010000100100";
		Trees_din <= x"009010a1";
		wait for Clk_period;
		Addr <=  "0010000100101";
		Trees_din <= x"17f77c04";
		wait for Clk_period;
		Addr <=  "0010000100110";
		Trees_din <= x"005d10a1";
		wait for Clk_period;
		Addr <=  "0010000100111";
		Trees_din <= x"ffcd10a1";
		wait for Clk_period;
		Addr <=  "0010000101000";
		Trees_din <= x"07fef114";
		wait for Clk_period;
		Addr <=  "0010000101001";
		Trees_din <= x"0005d210";
		wait for Clk_period;
		Addr <=  "0010000101010";
		Trees_din <= x"0003e304";
		wait for Clk_period;
		Addr <=  "0010000101011";
		Trees_din <= x"ff85116d";
		wait for Clk_period;
		Addr <=  "0010000101100";
		Trees_din <= x"08003f08";
		wait for Clk_period;
		Addr <=  "0010000101101";
		Trees_din <= x"0e002904";
		wait for Clk_period;
		Addr <=  "0010000101110";
		Trees_din <= x"ffb1116d";
		wait for Clk_period;
		Addr <=  "0010000101111";
		Trees_din <= x"00e9116d";
		wait for Clk_period;
		Addr <=  "0010000110000";
		Trees_din <= x"ffa2116d";
		wait for Clk_period;
		Addr <=  "0010000110001";
		Trees_din <= x"ff6b116d";
		wait for Clk_period;
		Addr <=  "0010000110010";
		Trees_din <= x"0703c32c";
		wait for Clk_period;
		Addr <=  "0010000110011";
		Trees_din <= x"00073710";
		wait for Clk_period;
		Addr <=  "0010000110100";
		Trees_din <= x"0a003b04";
		wait for Clk_period;
		Addr <=  "0010000110101";
		Trees_din <= x"0057116d";
		wait for Clk_period;
		Addr <=  "0010000110110";
		Trees_din <= x"010a8108";
		wait for Clk_period;
		Addr <=  "0010000110111";
		Trees_din <= x"010a6404";
		wait for Clk_period;
		Addr <=  "0010000111000";
		Trees_din <= x"ffc6116d";
		wait for Clk_period;
		Addr <=  "0010000111001";
		Trees_din <= x"00aa116d";
		wait for Clk_period;
		Addr <=  "0010000111010";
		Trees_din <= x"ff74116d";
		wait for Clk_period;
		Addr <=  "0010000111011";
		Trees_din <= x"12008310";
		wait for Clk_period;
		Addr <=  "0010000111100";
		Trees_din <= x"07030e08";
		wait for Clk_period;
		Addr <=  "0010000111101";
		Trees_din <= x"00080404";
		wait for Clk_period;
		Addr <=  "0010000111110";
		Trees_din <= x"0040116d";
		wait for Clk_period;
		Addr <=  "0010000111111";
		Trees_din <= x"ff7b116d";
		wait for Clk_period;
		Addr <=  "0010001000000";
		Trees_din <= x"11005c04";
		wait for Clk_period;
		Addr <=  "0010001000001";
		Trees_din <= x"008f116d";
		wait for Clk_period;
		Addr <=  "0010001000010";
		Trees_din <= x"0001116d";
		wait for Clk_period;
		Addr <=  "0010001000011";
		Trees_din <= x"0b008408";
		wait for Clk_period;
		Addr <=  "0010001000100";
		Trees_din <= x"06ff2a04";
		wait for Clk_period;
		Addr <=  "0010001000101";
		Trees_din <= x"013a116d";
		wait for Clk_period;
		Addr <=  "0010001000110";
		Trees_din <= x"0019116d";
		wait for Clk_period;
		Addr <=  "0010001000111";
		Trees_din <= x"ffea116d";
		wait for Clk_period;
		Addr <=  "0010001001000";
		Trees_din <= x"14021508";
		wait for Clk_period;
		Addr <=  "0010001001001";
		Trees_din <= x"0f00bc04";
		wait for Clk_period;
		Addr <=  "0010001001010";
		Trees_din <= x"0010116d";
		wait for Clk_period;
		Addr <=  "0010001001011";
		Trees_din <= x"ff85116d";
		wait for Clk_period;
		Addr <=  "0010001001100";
		Trees_din <= x"1800a210";
		wait for Clk_period;
		Addr <=  "0010001001101";
		Trees_din <= x"03f8ba08";
		wait for Clk_period;
		Addr <=  "0010001001110";
		Trees_din <= x"11001104";
		wait for Clk_period;
		Addr <=  "0010001001111";
		Trees_din <= x"0030116d";
		wait for Clk_period;
		Addr <=  "0010001010000";
		Trees_din <= x"ff97116d";
		wait for Clk_period;
		Addr <=  "0010001010001";
		Trees_din <= x"11010404";
		wait for Clk_period;
		Addr <=  "0010001010010";
		Trees_din <= x"004c116d";
		wait for Clk_period;
		Addr <=  "0010001010011";
		Trees_din <= x"ffd7116d";
		wait for Clk_period;
		Addr <=  "0010001010100";
		Trees_din <= x"04fab708";
		wait for Clk_period;
		Addr <=  "0010001010101";
		Trees_din <= x"1b028604";
		wait for Clk_period;
		Addr <=  "0010001010110";
		Trees_din <= x"ffd2116d";
		wait for Clk_period;
		Addr <=  "0010001010111";
		Trees_din <= x"0068116d";
		wait for Clk_period;
		Addr <=  "0010001011000";
		Trees_din <= x"00053f04";
		wait for Clk_period;
		Addr <=  "0010001011001";
		Trees_din <= x"008b116d";
		wait for Clk_period;
		Addr <=  "0010001011010";
		Trees_din <= x"fffc116d";
		wait for Clk_period;
		Addr <=  "0010001011011";
		Trees_din <= x"07fef114";
		wait for Clk_period;
		Addr <=  "0010001011100";
		Trees_din <= x"0005d210";
		wait for Clk_period;
		Addr <=  "0010001011101";
		Trees_din <= x"05f61a08";
		wait for Clk_period;
		Addr <=  "0010001011110";
		Trees_din <= x"05f56304";
		wait for Clk_period;
		Addr <=  "0010001011111";
		Trees_din <= x"ffa81219";
		wait for Clk_period;
		Addr <=  "0010001100000";
		Trees_din <= x"00d91219";
		wait for Clk_period;
		Addr <=  "0010001100001";
		Trees_din <= x"07fe6604";
		wait for Clk_period;
		Addr <=  "0010001100010";
		Trees_din <= x"ff841219";
		wait for Clk_period;
		Addr <=  "0010001100011";
		Trees_din <= x"00111219";
		wait for Clk_period;
		Addr <=  "0010001100100";
		Trees_din <= x"ff6c1219";
		wait for Clk_period;
		Addr <=  "0010001100101";
		Trees_din <= x"070c0a30";
		wait for Clk_period;
		Addr <=  "0010001100110";
		Trees_din <= x"0a003d18";
		wait for Clk_period;
		Addr <=  "0010001100111";
		Trees_din <= x"06fd7e08";
		wait for Clk_period;
		Addr <=  "0010001101000";
		Trees_din <= x"13037804";
		wait for Clk_period;
		Addr <=  "0010001101001";
		Trees_din <= x"fff41219";
		wait for Clk_period;
		Addr <=  "0010001101010";
		Trees_din <= x"ff8f1219";
		wait for Clk_period;
		Addr <=  "0010001101011";
		Trees_din <= x"04fd1d08";
		wait for Clk_period;
		Addr <=  "0010001101100";
		Trees_din <= x"11017504";
		wait for Clk_period;
		Addr <=  "0010001101101";
		Trees_din <= x"00db1219";
		wait for Clk_period;
		Addr <=  "0010001101110";
		Trees_din <= x"00191219";
		wait for Clk_period;
		Addr <=  "0010001101111";
		Trees_din <= x"19000f04";
		wait for Clk_period;
		Addr <=  "0010001110000";
		Trees_din <= x"ffa71219";
		wait for Clk_period;
		Addr <=  "0010001110001";
		Trees_din <= x"00381219";
		wait for Clk_period;
		Addr <=  "0010001110010";
		Trees_din <= x"07006c08";
		wait for Clk_period;
		Addr <=  "0010001110011";
		Trees_din <= x"1b024404";
		wait for Clk_period;
		Addr <=  "0010001110100";
		Trees_din <= x"00681219";
		wait for Clk_period;
		Addr <=  "0010001110101";
		Trees_din <= x"ff741219";
		wait for Clk_period;
		Addr <=  "0010001110110";
		Trees_din <= x"22000508";
		wait for Clk_period;
		Addr <=  "0010001110111";
		Trees_din <= x"0900f404";
		wait for Clk_period;
		Addr <=  "0010001111000";
		Trees_din <= x"00011219";
		wait for Clk_period;
		Addr <=  "0010001111001";
		Trees_din <= x"ff8b1219";
		wait for Clk_period;
		Addr <=  "0010001111010";
		Trees_din <= x"22000a04";
		wait for Clk_period;
		Addr <=  "0010001111011";
		Trees_din <= x"00b01219";
		wait for Clk_period;
		Addr <=  "0010001111100";
		Trees_din <= x"002f1219";
		wait for Clk_period;
		Addr <=  "0010001111101";
		Trees_din <= x"08003a08";
		wait for Clk_period;
		Addr <=  "0010001111110";
		Trees_din <= x"1c025104";
		wait for Clk_period;
		Addr <=  "0010001111111";
		Trees_din <= x"00561219";
		wait for Clk_period;
		Addr <=  "0010010000000";
		Trees_din <= x"ffb21219";
		wait for Clk_period;
		Addr <=  "0010010000001";
		Trees_din <= x"1303d404";
		wait for Clk_period;
		Addr <=  "0010010000010";
		Trees_din <= x"00891219";
		wait for Clk_period;
		Addr <=  "0010010000011";
		Trees_din <= x"17f77c04";
		wait for Clk_period;
		Addr <=  "0010010000100";
		Trees_din <= x"00561219";
		wait for Clk_period;
		Addr <=  "0010010000101";
		Trees_din <= x"ffd21219";
		wait for Clk_period;
		Addr <=  "0010010000110";
		Trees_din <= x"07fef114";
		wait for Clk_period;
		Addr <=  "0010010000111";
		Trees_din <= x"0005d210";
		wait for Clk_period;
		Addr <=  "0010010001000";
		Trees_din <= x"05f61a08";
		wait for Clk_period;
		Addr <=  "0010010001001";
		Trees_din <= x"05f56304";
		wait for Clk_period;
		Addr <=  "0010010001010";
		Trees_din <= x"ffac12bd";
		wait for Clk_period;
		Addr <=  "0010010001011";
		Trees_din <= x"00b712bd";
		wait for Clk_period;
		Addr <=  "0010010001100";
		Trees_din <= x"0401d104";
		wait for Clk_period;
		Addr <=  "0010010001101";
		Trees_din <= x"ff8912bd";
		wait for Clk_period;
		Addr <=  "0010010001110";
		Trees_din <= x"000a12bd";
		wait for Clk_period;
		Addr <=  "0010010001111";
		Trees_din <= x"ff6d12bd";
		wait for Clk_period;
		Addr <=  "0010010010000";
		Trees_din <= x"070c0a28";
		wait for Clk_period;
		Addr <=  "0010010010001";
		Trees_din <= x"02fe9208";
		wait for Clk_period;
		Addr <=  "0010010010010";
		Trees_din <= x"10003c04";
		wait for Clk_period;
		Addr <=  "0010010010011";
		Trees_din <= x"000e12bd";
		wait for Clk_period;
		Addr <=  "0010010010100";
		Trees_din <= x"ff7612bd";
		wait for Clk_period;
		Addr <=  "0010010010101";
		Trees_din <= x"05fb9610";
		wait for Clk_period;
		Addr <=  "0010010010110";
		Trees_din <= x"0b007808";
		wait for Clk_period;
		Addr <=  "0010010010111";
		Trees_din <= x"03fa3904";
		wait for Clk_period;
		Addr <=  "0010010011000";
		Trees_din <= x"ffac12bd";
		wait for Clk_period;
		Addr <=  "0010010011001";
		Trees_din <= x"001312bd";
		wait for Clk_period;
		Addr <=  "0010010011010";
		Trees_din <= x"06ff2a04";
		wait for Clk_period;
		Addr <=  "0010010011011";
		Trees_din <= x"004012bd";
		wait for Clk_period;
		Addr <=  "0010010011100";
		Trees_din <= x"ffda12bd";
		wait for Clk_period;
		Addr <=  "0010010011101";
		Trees_din <= x"05fdce08";
		wait for Clk_period;
		Addr <=  "0010010011110";
		Trees_din <= x"03f8ad04";
		wait for Clk_period;
		Addr <=  "0010010011111";
		Trees_din <= x"00ae12bd";
		wait for Clk_period;
		Addr <=  "0010010100000";
		Trees_din <= x"002c12bd";
		wait for Clk_period;
		Addr <=  "0010010100001";
		Trees_din <= x"1f025204";
		wait for Clk_period;
		Addr <=  "0010010100010";
		Trees_din <= x"006c12bd";
		wait for Clk_period;
		Addr <=  "0010010100011";
		Trees_din <= x"ffc612bd";
		wait for Clk_period;
		Addr <=  "0010010100100";
		Trees_din <= x"0f003710";
		wait for Clk_period;
		Addr <=  "0010010100101";
		Trees_din <= x"0f00050c";
		wait for Clk_period;
		Addr <=  "0010010100110";
		Trees_din <= x"010a6404";
		wait for Clk_period;
		Addr <=  "0010010100111";
		Trees_din <= x"006512bd";
		wait for Clk_period;
		Addr <=  "0010010101000";
		Trees_din <= x"0c008804";
		wait for Clk_period;
		Addr <=  "0010010101001";
		Trees_din <= x"000012bd";
		wait for Clk_period;
		Addr <=  "0010010101010";
		Trees_din <= x"ffcf12bd";
		wait for Clk_period;
		Addr <=  "0010010101011";
		Trees_din <= x"008612bd";
		wait for Clk_period;
		Addr <=  "0010010101100";
		Trees_din <= x"0c00a904";
		wait for Clk_period;
		Addr <=  "0010010101101";
		Trees_din <= x"001412bd";
		wait for Clk_period;
		Addr <=  "0010010101110";
		Trees_din <= x"ffd612bd";
		wait for Clk_period;
		Addr <=  "0010010101111";
		Trees_din <= x"07fef114";
		wait for Clk_period;
		Addr <=  "0010010110000";
		Trees_din <= x"0005d210";
		wait for Clk_period;
		Addr <=  "0010010110001";
		Trees_din <= x"0003e304";
		wait for Clk_period;
		Addr <=  "0010010110010";
		Trees_din <= x"ff8f1339";
		wait for Clk_period;
		Addr <=  "0010010110011";
		Trees_din <= x"0d005f04";
		wait for Clk_period;
		Addr <=  "0010010110100";
		Trees_din <= x"ffab1339";
		wait for Clk_period;
		Addr <=  "0010010110101";
		Trees_din <= x"0900d904";
		wait for Clk_period;
		Addr <=  "0010010110110";
		Trees_din <= x"fff81339";
		wait for Clk_period;
		Addr <=  "0010010110111";
		Trees_din <= x"00b21339";
		wait for Clk_period;
		Addr <=  "0010010111000";
		Trees_din <= x"ff6e1339";
		wait for Clk_period;
		Addr <=  "0010010111001";
		Trees_din <= x"1af94008";
		wait for Clk_period;
		Addr <=  "0010010111010";
		Trees_din <= x"0a004004";
		wait for Clk_period;
		Addr <=  "0010010111011";
		Trees_din <= x"00021339";
		wait for Clk_period;
		Addr <=  "0010010111100";
		Trees_din <= x"ff7e1339";
		wait for Clk_period;
		Addr <=  "0010010111101";
		Trees_din <= x"1300b208";
		wait for Clk_period;
		Addr <=  "0010010111110";
		Trees_din <= x"00ffa604";
		wait for Clk_period;
		Addr <=  "0010010111111";
		Trees_din <= x"ff801339";
		wait for Clk_period;
		Addr <=  "0010011000000";
		Trees_din <= x"ffe41339";
		wait for Clk_period;
		Addr <=  "0010011000001";
		Trees_din <= x"08004a10";
		wait for Clk_period;
		Addr <=  "0010011000010";
		Trees_din <= x"1e028508";
		wait for Clk_period;
		Addr <=  "0010011000011";
		Trees_din <= x"0900bd04";
		wait for Clk_period;
		Addr <=  "0010011000100";
		Trees_din <= x"ffd61339";
		wait for Clk_period;
		Addr <=  "0010011000101";
		Trees_din <= x"00121339";
		wait for Clk_period;
		Addr <=  "0010011000110";
		Trees_din <= x"0702a704";
		wait for Clk_period;
		Addr <=  "0010011000111";
		Trees_din <= x"ffc71339";
		wait for Clk_period;
		Addr <=  "0010011001000";
		Trees_din <= x"00771339";
		wait for Clk_period;
		Addr <=  "0010011001001";
		Trees_din <= x"1b026404";
		wait for Clk_period;
		Addr <=  "0010011001010";
		Trees_din <= x"ffc11339";
		wait for Clk_period;
		Addr <=  "0010011001011";
		Trees_din <= x"16006a04";
		wait for Clk_period;
		Addr <=  "0010011001100";
		Trees_din <= x"fff11339";
		wait for Clk_period;
		Addr <=  "0010011001101";
		Trees_din <= x"00851339";
		wait for Clk_period;
		Addr <=  "0010011001110";
		Trees_din <= x"07fe660c";
		wait for Clk_period;
		Addr <=  "0010011001111";
		Trees_din <= x"12005a04";
		wait for Clk_period;
		Addr <=  "0010011010000";
		Trees_din <= x"003513dd";
		wait for Clk_period;
		Addr <=  "0010011010001";
		Trees_din <= x"1d028604";
		wait for Clk_period;
		Addr <=  "0010011010010";
		Trees_din <= x"ff6e13dd";
		wait for Clk_period;
		Addr <=  "0010011010011";
		Trees_din <= x"001f13dd";
		wait for Clk_period;
		Addr <=  "0010011010100";
		Trees_din <= x"0207fb40";
		wait for Clk_period;
		Addr <=  "0010011010101";
		Trees_din <= x"10004620";
		wait for Clk_period;
		Addr <=  "0010011010110";
		Trees_din <= x"04fc9610";
		wait for Clk_period;
		Addr <=  "0010011010111";
		Trees_din <= x"16006a08";
		wait for Clk_period;
		Addr <=  "0010011011000";
		Trees_din <= x"18010c04";
		wait for Clk_period;
		Addr <=  "0010011011001";
		Trees_din <= x"004f13dd";
		wait for Clk_period;
		Addr <=  "0010011011010";
		Trees_din <= x"ffd813dd";
		wait for Clk_period;
		Addr <=  "0010011011011";
		Trees_din <= x"12007104";
		wait for Clk_period;
		Addr <=  "0010011011100";
		Trees_din <= x"002513dd";
		wait for Clk_period;
		Addr <=  "0010011011101";
		Trees_din <= x"ff7813dd";
		wait for Clk_period;
		Addr <=  "0010011011110";
		Trees_din <= x"0d017008";
		wait for Clk_period;
		Addr <=  "0010011011111";
		Trees_din <= x"16004f04";
		wait for Clk_period;
		Addr <=  "0010011100000";
		Trees_din <= x"ffff13dd";
		wait for Clk_period;
		Addr <=  "0010011100001";
		Trees_din <= x"ff6c13dd";
		wait for Clk_period;
		Addr <=  "0010011100010";
		Trees_din <= x"04fd8b04";
		wait for Clk_period;
		Addr <=  "0010011100011";
		Trees_din <= x"ffb613dd";
		wait for Clk_period;
		Addr <=  "0010011100100";
		Trees_din <= x"007d13dd";
		wait for Clk_period;
		Addr <=  "0010011100101";
		Trees_din <= x"01063110";
		wait for Clk_period;
		Addr <=  "0010011100110";
		Trees_din <= x"0a005408";
		wait for Clk_period;
		Addr <=  "0010011100111";
		Trees_din <= x"07030e04";
		wait for Clk_period;
		Addr <=  "0010011101000";
		Trees_din <= x"000a13dd";
		wait for Clk_period;
		Addr <=  "0010011101001";
		Trees_din <= x"008b13dd";
		wait for Clk_period;
		Addr <=  "0010011101010";
		Trees_din <= x"02043b04";
		wait for Clk_period;
		Addr <=  "0010011101011";
		Trees_din <= x"002113dd";
		wait for Clk_period;
		Addr <=  "0010011101100";
		Trees_din <= x"ff9d13dd";
		wait for Clk_period;
		Addr <=  "0010011101101";
		Trees_din <= x"05f98208";
		wait for Clk_period;
		Addr <=  "0010011101110";
		Trees_din <= x"16007304";
		wait for Clk_period;
		Addr <=  "0010011101111";
		Trees_din <= x"005b13dd";
		wait for Clk_period;
		Addr <=  "0010011110000";
		Trees_din <= x"fffa13dd";
		wait for Clk_period;
		Addr <=  "0010011110001";
		Trees_din <= x"0c009304";
		wait for Clk_period;
		Addr <=  "0010011110010";
		Trees_din <= x"001e13dd";
		wait for Clk_period;
		Addr <=  "0010011110011";
		Trees_din <= x"ff6513dd";
		wait for Clk_period;
		Addr <=  "0010011110100";
		Trees_din <= x"0602d004";
		wait for Clk_period;
		Addr <=  "0010011110101";
		Trees_din <= x"ff8213dd";
		wait for Clk_period;
		Addr <=  "0010011110110";
		Trees_din <= x"002a13dd";
		wait for Clk_period;
		Addr <=  "0010011110111";
		Trees_din <= x"07fe660c";
		wait for Clk_period;
		Addr <=  "0010011111000";
		Trees_din <= x"0005d208";
		wait for Clk_period;
		Addr <=  "0010011111001";
		Trees_din <= x"05f61a04";
		wait for Clk_period;
		Addr <=  "0010011111010";
		Trees_din <= x"005514a1";
		wait for Clk_period;
		Addr <=  "0010011111011";
		Trees_din <= x"ff9314a1";
		wait for Clk_period;
		Addr <=  "0010011111100";
		Trees_din <= x"ff7114a1";
		wait for Clk_period;
		Addr <=  "0010011111101";
		Trees_din <= x"07047420";
		wait for Clk_period;
		Addr <=  "0010011111110";
		Trees_din <= x"02021704";
		wait for Clk_period;
		Addr <=  "0010011111111";
		Trees_din <= x"ff7714a1";
		wait for Clk_period;
		Addr <=  "0010100000000";
		Trees_din <= x"0204d90c";
		wait for Clk_period;
		Addr <=  "0010100000001";
		Trees_din <= x"10003e04";
		wait for Clk_period;
		Addr <=  "0010100000010";
		Trees_din <= x"ff9614a1";
		wait for Clk_period;
		Addr <=  "0010100000011";
		Trees_din <= x"010e3204";
		wait for Clk_period;
		Addr <=  "0010100000100";
		Trees_din <= x"005c14a1";
		wait for Clk_period;
		Addr <=  "0010100000101";
		Trees_din <= x"ffc514a1";
		wait for Clk_period;
		Addr <=  "0010100000110";
		Trees_din <= x"0900ef08";
		wait for Clk_period;
		Addr <=  "0010100000111";
		Trees_din <= x"19000304";
		wait for Clk_period;
		Addr <=  "0010100001000";
		Trees_din <= x"ff8314a1";
		wait for Clk_period;
		Addr <=  "0010100001001";
		Trees_din <= x"002114a1";
		wait for Clk_period;
		Addr <=  "0010100001010";
		Trees_din <= x"1303e804";
		wait for Clk_period;
		Addr <=  "0010100001011";
		Trees_din <= x"ffa714a1";
		wait for Clk_period;
		Addr <=  "0010100001100";
		Trees_din <= x"007714a1";
		wait for Clk_period;
		Addr <=  "0010100001101";
		Trees_din <= x"0900e720";
		wait for Clk_period;
		Addr <=  "0010100001110";
		Trees_din <= x"0900b810";
		wait for Clk_period;
		Addr <=  "0010100001111";
		Trees_din <= x"0706bc08";
		wait for Clk_period;
		Addr <=  "0010100010000";
		Trees_din <= x"04fccc04";
		wait for Clk_period;
		Addr <=  "0010100010001";
		Trees_din <= x"ff8214a1";
		wait for Clk_period;
		Addr <=  "0010100010010";
		Trees_din <= x"002214a1";
		wait for Clk_period;
		Addr <=  "0010100010011";
		Trees_din <= x"04faec04";
		wait for Clk_period;
		Addr <=  "0010100010100";
		Trees_din <= x"ffee14a1";
		wait for Clk_period;
		Addr <=  "0010100010101";
		Trees_din <= x"006414a1";
		wait for Clk_period;
		Addr <=  "0010100010110";
		Trees_din <= x"03f7e708";
		wait for Clk_period;
		Addr <=  "0010100010111";
		Trees_din <= x"02023a04";
		wait for Clk_period;
		Addr <=  "0010100011000";
		Trees_din <= x"005714a1";
		wait for Clk_period;
		Addr <=  "0010100011001";
		Trees_din <= x"ff9c14a1";
		wait for Clk_period;
		Addr <=  "0010100011010";
		Trees_din <= x"0f007f04";
		wait for Clk_period;
		Addr <=  "0010100011011";
		Trees_din <= x"008d14a1";
		wait for Clk_period;
		Addr <=  "0010100011100";
		Trees_din <= x"fffc14a1";
		wait for Clk_period;
		Addr <=  "0010100011101";
		Trees_din <= x"10004710";
		wait for Clk_period;
		Addr <=  "0010100011110";
		Trees_din <= x"05fa8508";
		wait for Clk_period;
		Addr <=  "0010100011111";
		Trees_din <= x"05f65604";
		wait for Clk_period;
		Addr <=  "0010100100000";
		Trees_din <= x"ffee14a1";
		wait for Clk_period;
		Addr <=  "0010100100001";
		Trees_din <= x"ff5514a1";
		wait for Clk_period;
		Addr <=  "0010100100010";
		Trees_din <= x"04fbee04";
		wait for Clk_period;
		Addr <=  "0010100100011";
		Trees_din <= x"006014a1";
		wait for Clk_period;
		Addr <=  "0010100100100";
		Trees_din <= x"ffc314a1";
		wait for Clk_period;
		Addr <=  "0010100100101";
		Trees_din <= x"04fa9604";
		wait for Clk_period;
		Addr <=  "0010100100110";
		Trees_din <= x"ffce14a1";
		wait for Clk_period;
		Addr <=  "0010100100111";
		Trees_din <= x"007614a1";
		wait for Clk_period;
		Addr <=  "0010100101000";
		Trees_din <= x"07fbbc04";
		wait for Clk_period;
		Addr <=  "0010100101001";
		Trees_din <= x"ff75153d";
		wait for Clk_period;
		Addr <=  "0010100101010";
		Trees_din <= x"07047420";
		wait for Clk_period;
		Addr <=  "0010100101011";
		Trees_din <= x"02021704";
		wait for Clk_period;
		Addr <=  "0010100101100";
		Trees_din <= x"ff7a153d";
		wait for Clk_period;
		Addr <=  "0010100101101";
		Trees_din <= x"0900ef10";
		wait for Clk_period;
		Addr <=  "0010100101110";
		Trees_din <= x"0900dd08";
		wait for Clk_period;
		Addr <=  "0010100101111";
		Trees_din <= x"0f000404";
		wait for Clk_period;
		Addr <=  "0010100110000";
		Trees_din <= x"ff8b153d";
		wait for Clk_period;
		Addr <=  "0010100110001";
		Trees_din <= x"0021153d";
		wait for Clk_period;
		Addr <=  "0010100110010";
		Trees_din <= x"0f000204";
		wait for Clk_period;
		Addr <=  "0010100110011";
		Trees_din <= x"001d153d";
		wait for Clk_period;
		Addr <=  "0010100110100";
		Trees_din <= x"ff75153d";
		wait for Clk_period;
		Addr <=  "0010100110101";
		Trees_din <= x"0d000004";
		wait for Clk_period;
		Addr <=  "0010100110110";
		Trees_din <= x"ffaa153d";
		wait for Clk_period;
		Addr <=  "0010100110111";
		Trees_din <= x"1100fe04";
		wait for Clk_period;
		Addr <=  "0010100111000";
		Trees_din <= x"0085153d";
		wait for Clk_period;
		Addr <=  "0010100111001";
		Trees_din <= x"ffe2153d";
		wait for Clk_period;
		Addr <=  "0010100111010";
		Trees_din <= x"0900e718";
		wait for Clk_period;
		Addr <=  "0010100111011";
		Trees_din <= x"17f72208";
		wait for Clk_period;
		Addr <=  "0010100111100";
		Trees_din <= x"00ffa604";
		wait for Clk_period;
		Addr <=  "0010100111101";
		Trees_din <= x"ffea153d";
		wait for Clk_period;
		Addr <=  "0010100111110";
		Trees_din <= x"00a9153d";
		wait for Clk_period;
		Addr <=  "0010100111111";
		Trees_din <= x"03f8f508";
		wait for Clk_period;
		Addr <=  "0010101000000";
		Trees_din <= x"0d00aa04";
		wait for Clk_period;
		Addr <=  "0010101000001";
		Trees_din <= x"ffa6153d";
		wait for Clk_period;
		Addr <=  "0010101000010";
		Trees_din <= x"001e153d";
		wait for Clk_period;
		Addr <=  "0010101000011";
		Trees_din <= x"02064e04";
		wait for Clk_period;
		Addr <=  "0010101000100";
		Trees_din <= x"0039153d";
		wait for Clk_period;
		Addr <=  "0010101000101";
		Trees_din <= x"ff8c153d";
		wait for Clk_period;
		Addr <=  "0010101000110";
		Trees_din <= x"01084c08";
		wait for Clk_period;
		Addr <=  "0010101000111";
		Trees_din <= x"06ff8e04";
		wait for Clk_period;
		Addr <=  "0010101001000";
		Trees_din <= x"0067153d";
		wait for Clk_period;
		Addr <=  "0010101001001";
		Trees_din <= x"ffc9153d";
		wait for Clk_period;
		Addr <=  "0010101001010";
		Trees_din <= x"05f5b004";
		wait for Clk_period;
		Addr <=  "0010101001011";
		Trees_din <= x"0037153d";
		wait for Clk_period;
		Addr <=  "0010101001100";
		Trees_din <= x"03f8d104";
		wait for Clk_period;
		Addr <=  "0010101001101";
		Trees_din <= x"ffd3153d";
		wait for Clk_period;
		Addr <=  "0010101001110";
		Trees_din <= x"ff48153d";
		wait for Clk_period;
		Addr <=  "0010101001111";
		Trees_din <= x"07fbbc04";
		wait for Clk_period;
		Addr <=  "0010101010000";
		Trees_din <= x"ff7715f9";
		wait for Clk_period;
		Addr <=  "0010101010001";
		Trees_din <= x"0204d93c";
		wait for Clk_period;
		Addr <=  "0010101010010";
		Trees_din <= x"1f026520";
		wait for Clk_period;
		Addr <=  "0010101010011";
		Trees_din <= x"0d003210";
		wait for Clk_period;
		Addr <=  "0010101010100";
		Trees_din <= x"1e025b08";
		wait for Clk_period;
		Addr <=  "0010101010101";
		Trees_din <= x"0c009d04";
		wait for Clk_period;
		Addr <=  "0010101010110";
		Trees_din <= x"002f15f9";
		wait for Clk_period;
		Addr <=  "0010101010111";
		Trees_din <= x"ff8415f9";
		wait for Clk_period;
		Addr <=  "0010101011000";
		Trees_din <= x"06fe6604";
		wait for Clk_period;
		Addr <=  "0010101011001";
		Trees_din <= x"007f15f9";
		wait for Clk_period;
		Addr <=  "0010101011010";
		Trees_din <= x"ffdf15f9";
		wait for Clk_period;
		Addr <=  "0010101011011";
		Trees_din <= x"04fad708";
		wait for Clk_period;
		Addr <=  "0010101011100";
		Trees_din <= x"0f000704";
		wait for Clk_period;
		Addr <=  "0010101011101";
		Trees_din <= x"ff9e15f9";
		wait for Clk_period;
		Addr <=  "0010101011110";
		Trees_din <= x"002515f9";
		wait for Clk_period;
		Addr <=  "0010101011111";
		Trees_din <= x"0005b004";
		wait for Clk_period;
		Addr <=  "0010101100000";
		Trees_din <= x"00b315f9";
		wait for Clk_period;
		Addr <=  "0010101100001";
		Trees_din <= x"001e15f9";
		wait for Clk_period;
		Addr <=  "0010101100010";
		Trees_din <= x"1afc1310";
		wait for Clk_period;
		Addr <=  "0010101100011";
		Trees_din <= x"0f002d08";
		wait for Clk_period;
		Addr <=  "0010101100100";
		Trees_din <= x"0b006804";
		wait for Clk_period;
		Addr <=  "0010101100101";
		Trees_din <= x"ffa915f9";
		wait for Clk_period;
		Addr <=  "0010101100110";
		Trees_din <= x"005515f9";
		wait for Clk_period;
		Addr <=  "0010101100111";
		Trees_din <= x"1f028604";
		wait for Clk_period;
		Addr <=  "0010101101000";
		Trees_din <= x"ffc315f9";
		wait for Clk_period;
		Addr <=  "0010101101001";
		Trees_din <= x"004715f9";
		wait for Clk_period;
		Addr <=  "0010101101010";
		Trees_din <= x"0f000808";
		wait for Clk_period;
		Addr <=  "0010101101011";
		Trees_din <= x"0109a704";
		wait for Clk_period;
		Addr <=  "0010101101100";
		Trees_din <= x"004f15f9";
		wait for Clk_period;
		Addr <=  "0010101101101";
		Trees_din <= x"ffaa15f9";
		wait for Clk_period;
		Addr <=  "0010101101110";
		Trees_din <= x"ff7e15f9";
		wait for Clk_period;
		Addr <=  "0010101101111";
		Trees_din <= x"0f000204";
		wait for Clk_period;
		Addr <=  "0010101110000";
		Trees_din <= x"ff7b15f9";
		wait for Clk_period;
		Addr <=  "0010101110001";
		Trees_din <= x"01026d0c";
		wait for Clk_period;
		Addr <=  "0010101110010";
		Trees_din <= x"06ff0804";
		wait for Clk_period;
		Addr <=  "0010101110011";
		Trees_din <= x"ff9b15f9";
		wait for Clk_period;
		Addr <=  "0010101110100";
		Trees_din <= x"04fe0c04";
		wait for Clk_period;
		Addr <=  "0010101110101";
		Trees_din <= x"000215f9";
		wait for Clk_period;
		Addr <=  "0010101110110";
		Trees_din <= x"009e15f9";
		wait for Clk_period;
		Addr <=  "0010101110111";
		Trees_din <= x"04fd1d08";
		wait for Clk_period;
		Addr <=  "0010101111000";
		Trees_din <= x"05f70f04";
		wait for Clk_period;
		Addr <=  "0010101111001";
		Trees_din <= x"002615f9";
		wait for Clk_period;
		Addr <=  "0010101111010";
		Trees_din <= x"ff9015f9";
		wait for Clk_period;
		Addr <=  "0010101111011";
		Trees_din <= x"18020204";
		wait for Clk_period;
		Addr <=  "0010101111100";
		Trees_din <= x"ff7815f9";
		wait for Clk_period;
		Addr <=  "0010101111101";
		Trees_din <= x"ffd515f9";
		wait for Clk_period;
		Addr <=  "0010101111110";
		Trees_din <= x"07fbbc04";
		wait for Clk_period;
		Addr <=  "0010101111111";
		Trees_din <= x"ff7a1685";
		wait for Clk_period;
		Addr <=  "0010110000000";
		Trees_din <= x"070d1338";
		wait for Clk_period;
		Addr <=  "0010110000001";
		Trees_din <= x"06fdee18";
		wait for Clk_period;
		Addr <=  "0010110000010";
		Trees_din <= x"06fc5f0c";
		wait for Clk_period;
		Addr <=  "0010110000011";
		Trees_din <= x"0f00bc08";
		wait for Clk_period;
		Addr <=  "0010110000100";
		Trees_din <= x"06fa9004";
		wait for Clk_period;
		Addr <=  "0010110000101";
		Trees_din <= x"ffda1685";
		wait for Clk_period;
		Addr <=  "0010110000110";
		Trees_din <= x"00411685";
		wait for Clk_period;
		Addr <=  "0010110000111";
		Trees_din <= x"ff851685";
		wait for Clk_period;
		Addr <=  "0010110001000";
		Trees_din <= x"0a005608";
		wait for Clk_period;
		Addr <=  "0010110001001";
		Trees_din <= x"07076704";
		wait for Clk_period;
		Addr <=  "0010110001010";
		Trees_din <= x"ff6d1685";
		wait for Clk_period;
		Addr <=  "0010110001011";
		Trees_din <= x"ffdd1685";
		wait for Clk_period;
		Addr <=  "0010110001100";
		Trees_din <= x"00411685";
		wait for Clk_period;
		Addr <=  "0010110001101";
		Trees_din <= x"06ff3110";
		wait for Clk_period;
		Addr <=  "0010110001110";
		Trees_din <= x"0c00ad08";
		wait for Clk_period;
		Addr <=  "0010110001111";
		Trees_din <= x"03fc5c04";
		wait for Clk_period;
		Addr <=  "0010110010000";
		Trees_din <= x"ffcb1685";
		wait for Clk_period;
		Addr <=  "0010110010001";
		Trees_din <= x"00811685";
		wait for Clk_period;
		Addr <=  "0010110010010";
		Trees_din <= x"08003804";
		wait for Clk_period;
		Addr <=  "0010110010011";
		Trees_din <= x"00231685";
		wait for Clk_period;
		Addr <=  "0010110010100";
		Trees_din <= x"009c1685";
		wait for Clk_period;
		Addr <=  "0010110010101";
		Trees_din <= x"01036908";
		wait for Clk_period;
		Addr <=  "0010110010110";
		Trees_din <= x"0e002904";
		wait for Clk_period;
		Addr <=  "0010110010111";
		Trees_din <= x"ffc51685";
		wait for Clk_period;
		Addr <=  "0010110011000";
		Trees_din <= x"00521685";
		wait for Clk_period;
		Addr <=  "0010110011001";
		Trees_din <= x"0d00ed04";
		wait for Clk_period;
		Addr <=  "0010110011010";
		Trees_din <= x"ffaa1685";
		wait for Clk_period;
		Addr <=  "0010110011011";
		Trees_din <= x"00091685";
		wait for Clk_period;
		Addr <=  "0010110011100";
		Trees_din <= x"18003108";
		wait for Clk_period;
		Addr <=  "0010110011101";
		Trees_din <= x"05f77a04";
		wait for Clk_period;
		Addr <=  "0010110011110";
		Trees_din <= x"ffcc1685";
		wait for Clk_period;
		Addr <=  "0010110011111";
		Trees_din <= x"002e1685";
		wait for Clk_period;
		Addr <=  "0010110100000";
		Trees_din <= x"00741685";
		wait for Clk_period;
		Addr <=  "0010110100001";
		Trees_din <= x"07fbbc04";
		wait for Clk_period;
		Addr <=  "0010110100010";
		Trees_din <= x"ff7c1721";
		wait for Clk_period;
		Addr <=  "0010110100011";
		Trees_din <= x"0b00631c";
		wait for Clk_period;
		Addr <=  "0010110100100";
		Trees_din <= x"04fd1d14";
		wait for Clk_period;
		Addr <=  "0010110100101";
		Trees_din <= x"0e004d10";
		wait for Clk_period;
		Addr <=  "0010110100110";
		Trees_din <= x"0204f408";
		wait for Clk_period;
		Addr <=  "0010110100111";
		Trees_din <= x"1b027c04";
		wait for Clk_period;
		Addr <=  "0010110101000";
		Trees_din <= x"008e1721";
		wait for Clk_period;
		Addr <=  "0010110101001";
		Trees_din <= x"001b1721";
		wait for Clk_period;
		Addr <=  "0010110101010";
		Trees_din <= x"10004a04";
		wait for Clk_period;
		Addr <=  "0010110101011";
		Trees_din <= x"003c1721";
		wait for Clk_period;
		Addr <=  "0010110101100";
		Trees_din <= x"ffc31721";
		wait for Clk_period;
		Addr <=  "0010110101101";
		Trees_din <= x"ffe01721";
		wait for Clk_period;
		Addr <=  "0010110101110";
		Trees_din <= x"0e004004";
		wait for Clk_period;
		Addr <=  "0010110101111";
		Trees_din <= x"00091721";
		wait for Clk_period;
		Addr <=  "0010110110000";
		Trees_din <= x"ff9a1721";
		wait for Clk_period;
		Addr <=  "0010110110001";
		Trees_din <= x"0b006814";
		wait for Clk_period;
		Addr <=  "0010110110010";
		Trees_din <= x"12006f08";
		wait for Clk_period;
		Addr <=  "0010110110011";
		Trees_din <= x"08004304";
		wait for Clk_period;
		Addr <=  "0010110110100";
		Trees_din <= x"ffbe1721";
		wait for Clk_period;
		Addr <=  "0010110110101";
		Trees_din <= x"00551721";
		wait for Clk_period;
		Addr <=  "0010110110110";
		Trees_din <= x"10004404";
		wait for Clk_period;
		Addr <=  "0010110110111";
		Trees_din <= x"fff91721";
		wait for Clk_period;
		Addr <=  "0010110111000";
		Trees_din <= x"05fb3104";
		wait for Clk_period;
		Addr <=  "0010110111001";
		Trees_din <= x"ff6d1721";
		wait for Clk_period;
		Addr <=  "0010110111010";
		Trees_din <= x"ffd21721";
		wait for Clk_period;
		Addr <=  "0010110111011";
		Trees_din <= x"07021b0c";
		wait for Clk_period;
		Addr <=  "0010110111100";
		Trees_din <= x"18015108";
		wait for Clk_period;
		Addr <=  "0010110111101";
		Trees_din <= x"1403d204";
		wait for Clk_period;
		Addr <=  "0010110111110";
		Trees_din <= x"008c1721";
		wait for Clk_period;
		Addr <=  "0010110111111";
		Trees_din <= x"ffd41721";
		wait for Clk_period;
		Addr <=  "0010111000000";
		Trees_din <= x"ff7e1721";
		wait for Clk_period;
		Addr <=  "0010111000001";
		Trees_din <= x"11014308";
		wait for Clk_period;
		Addr <=  "0010111000010";
		Trees_din <= x"1303df04";
		wait for Clk_period;
		Addr <=  "0010111000011";
		Trees_din <= x"ffa21721";
		wait for Clk_period;
		Addr <=  "0010111000100";
		Trees_din <= x"00151721";
		wait for Clk_period;
		Addr <=  "0010111000101";
		Trees_din <= x"19000a04";
		wait for Clk_period;
		Addr <=  "0010111000110";
		Trees_din <= x"00101721";
		wait for Clk_period;
		Addr <=  "0010111000111";
		Trees_din <= x"00691721";
		wait for Clk_period;
		Addr <=  "0010111001000";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  3
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"0307c234";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"0300dc18";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"03fee00c";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"0a005f04";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"ff5100a5";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"02070c04";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"ff8100a5";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"003700a5";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"17faaa08";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"1afd8b04";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"ff5c00a5";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"003700a5";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"00c200a5";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"04f92e08";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"00036a04";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"ff5f00a5";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"002100a5";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"10005610";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"0f000708";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"0a004604";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"ff7300a5";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"003700a5";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"0f001704";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"018d00a5";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"ffde00a5";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"023500a5";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"030e8418";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"04f77008";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"01091704";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"003700a5";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"ff9c00a5";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"02087008";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"06f8d704";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"00df00a5";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"039100a5";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"00000e04";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"ffa400a5";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"00ca00a5";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"1cfec804";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"015c00a5";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"048700a5";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"0305a72c";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"03fee00c";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"1d028804";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"ff570141";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"0d000904";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"003f0141";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"ff910141";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"04fa4308";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"0900ec04";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"ff5f0141";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"fff70141";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"0c00a60c";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"03033e08";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"0d003904";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"ffb00141";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"01000141";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"01c30141";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"1d024104";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"00760141";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"19001204";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"ff650141";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"00270141";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"010e8420";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"01079710";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"0e001004";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"00240141";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"0c005e04";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"00670141";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"14011a04";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"00c10141";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"01bb0141";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"0208530c";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"0a004d08";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"02027604";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"00090141";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"017a0141";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"fff90141";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"ff9f0141";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"ff960141";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"03045c2c";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"03fee00c";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"1f052404";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"ff5a01e5";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"18013304";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"ff9701e5";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"003f01e5";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"0203bf04";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"ff6201e5";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"0204d90c";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"0b007408";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"0900d104";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"006501e5";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"022301e5";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"ff9e01e5";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"09008108";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"09006e04";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"ff9f01e5";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"011701e5";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"0a004904";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"ff6901e5";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"001c01e5";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"030c2c18";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"05f56804";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"ff7201e5";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"00fcf308";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"0b006d04";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"ff7f01e5";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"002a01e5";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"0d01e808";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"0f001404";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"016e01e5";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"009101e5";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"ff9c01e5";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"010c730c";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"08004d08";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"1cfec804";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"005a01e5";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"013701e5";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"006701e5";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"005701e5";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"03045c34";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"03fee014";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"1d02880c";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"03fca204";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"ff5c02b1";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"0b009904";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"ff6402b1";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"009a02b1";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"05f64604";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"ffa402b1";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"004302b1";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"0203bf04";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"ff6702b1";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"0204d90c";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"0b007408";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"0900d104";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"005802b1";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"019d02b1";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"ffa602b1";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"09008108";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"09006e04";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"ffa402b1";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"00ee02b1";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"0a004904";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"ff6e02b1";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"001c02b1";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"030c2c1c";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"05f56804";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"ff7902b1";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"00fcf308";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"05f89e04";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"002102b1";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"ff8102b1";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"0b006408";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"06fb7504";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"ff7c02b1";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"00b602b1";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"0c00b204";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"011b02b1";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"003202b1";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"04f60108";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"030e8404";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"ffa502b1";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"00b802b1";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"1ff9f804";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"005002b1";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"11000004";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"004502b1";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"0a005604";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"00fd02b1";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"007802b1";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"03033e28";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"03fee010";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"0a005f0c";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"03fca204";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"ff5e036d";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"0b009904";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"ff68036d";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"008d036d";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"fffc036d";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"0203bf04";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"ff6f036d";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"0204d90c";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"0900d308";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"00025504";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"ffa1036d";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"00a2036d";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"011a036d";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"1e028704";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"ff6e036d";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"008f036d";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"030c2c1c";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"05f57104";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"ff7a036d";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"00fcf308";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"010ab104";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"ff74036d";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"0027036d";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"07027d08";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"0a003d04";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"fff5036d";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"0106036d";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"08003b04";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"ff64036d";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"008d036d";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"0700f908";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"1cfec804";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"0043036d";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"00e1036d";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"0d000308";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"05f62204";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"ff80036d";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"0041036d";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"0701a008";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"0a004804";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"0088036d";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"ff45036d";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"00f3036d";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"03033e28";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"03fee010";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"1f05240c";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"03fca204";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"ff600431";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"0e001d04";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"008a0431";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"ff6b0431";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"00040431";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"0203bf04";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"ff740431";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"0204d90c";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"0900d308";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"0c009504";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"ffa00431";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"009b0431";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"00f10431";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"1e028704";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"ff720431";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"00840431";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"030c2c1c";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"05f57104";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"ff800431";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"00fcf308";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"02037504";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"001a0431";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"ff790431";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"07027d08";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"0a003d04";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"fff30431";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"00d60431";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"08003b04";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"ff6b0431";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"00700431";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"0700f908";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"1cfec804";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"00350431";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"00ca0431";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"0d000308";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"05f62204";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"ff860431";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"00350431";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"0701a008";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"0a004804";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"00700431";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"ff550431";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"14021504";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"003d0431";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"00e20431";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"03033e28";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"03fee010";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"1d02880c";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"03fca204";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"ff6104dd";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"08003004";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"007c04dd";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"ff6e04dd";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"001604dd";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"04fb0208";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"1afa6704";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"003004dd";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"ff7304dd";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"01049404";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"ff8d04dd";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"010e6308";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"0204d904";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"00e104dd";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"001804dd";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"ffa504dd";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"0700f910";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"1cfec804";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"002704dd";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"0307c208";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"08003d04";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"00ab04dd";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"ff9a04dd";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"00ba04dd";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"03103e18";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"0205c80c";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"010e8408";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"01001d04";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"ffbf04dd";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"009604dd";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"ff9c04dd";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"06fc8b08";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"05f62b04";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"001b04dd";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"ff6304dd";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"00ad04dd";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"07012a04";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"ffee04dd";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"00bc04dd";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"0300dc24";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"03fdcb10";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"0a005f0c";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"0e001208";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"1d027404";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"ff9205a9";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"004505a9";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"ff6205a9";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"002305a9";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"1802330c";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"010d9f04";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"ff7305a9";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"010e6304";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"00aa05a9";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"ff9205a9";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"08004004";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"011605a9";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"ffae05a9";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"030c2c24";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"06f9bc10";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"0106ed08";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"01064904";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"ffd905a9";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"009205a9";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"08004504";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"ff6f05a9";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"ffe505a9";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"10005610";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"12006f08";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"0203d804";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"000d05a9";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"ff7505a9";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"0c00ac04";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"008c05a9";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"fff105a9";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"00d505a9";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"1ff9f804";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"fff205a9";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"0700f90c";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"1efd9f04";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"002305a9";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"020b5c04";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"00b705a9";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"006605a9";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"0701a008";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"01046504";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"009305a9";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"ff9f05a9";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"0d000304";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"ff9105a9";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"00c605a9";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"03fee010";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"1f05240c";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"03fca204";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"ff630649";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"0b009904";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"ff760649";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"00830649";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"002b0649";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"030c2c1c";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"1af96708";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"1801d904";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"00c30649";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"00290649";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"1f027b0c";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"00fd1a04";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"ff710649";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"05f43904";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"ff8d0649";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"00450649";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"1af9e504";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"00030649";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"ff650649";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"19000114";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"020b5c0c";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"0b009404";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"00b50649";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"02083e04";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"ffc50649";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"006b0649";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"0b006a04";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"ff9a0649";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"008b0649";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"03145b0c";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"19000304";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"ff5b0649";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"020a1604";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"00910649";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"ffb00649";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"00a60649";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"03fee010";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"0a005f0c";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"03fca204";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"ff6406dd";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"0e001d04";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"007406dd";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"ff7906dd";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"003506dd";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"030c2c1c";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"10005614";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"1af8eb04";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"00a106dd";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"0b006808";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"00078204";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"ff6306dd";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"006f06dd";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"12007704";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"006106dd";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"ffc706dd";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"10005c04";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"00ca06dd";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"fff006dd";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"19000110";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"020b5c08";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"0b009404";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"00ad06dd";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"001606dd";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"0b006a04";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"ffa106dd";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"008106dd";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"03145b0c";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"19000304";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"ff6706dd";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"020a1604";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"008806dd";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"ffb606dd";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"009d06dd";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"03fee010";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"1d02880c";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"03fca204";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"ff650789";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"0b009904";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"ff7d0789";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"00650789";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"003e0789";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"03103e34";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"17f76914";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"0704a90c";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"08003604";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"ffde0789";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"06fc5604";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"00c40789";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"001f0789";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"0b006804";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"ffa90789";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"00020789";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"1303ad10";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"19000708";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"17f82404";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"003c0789";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"ff6f0789";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"09007804";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"000e0789";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"00b50789";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"15003108";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"0107ec04";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"00880789";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"ffeb0789";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"0f000804";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"00090789";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"ff6f0789";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"020b5c0c";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"010a9f08";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"0001a204";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"00a50789";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"00090789";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"000b0789";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"04f97604";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"007a0789";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"ff9c0789";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"03fee010";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"1f05240c";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"03fca204";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"ff650835";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"08003004";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"005f0835";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"ff810835";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"00400835";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"030c2c24";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"1000561c";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"0c00970c";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"00059d08";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"08003404";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"ffef0835";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"ff6c0835";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"005c0835";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"0c00b208";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"04f91b04";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"ffe90835";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"00620835";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"04fce804";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"ff9a0835";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"00970835";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"10005c04";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"00ac0835";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"fff20835";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"19000114";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"020b5c0c";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"0b008e04";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"00a70835";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"07013e04";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"006b0835";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"ffb60835";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"0b006a04";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"ff9d0835";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"00760835";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"03145b0c";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"19000304";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"ff780835";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"020a1604";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"007b0835";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"ffc30835";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"00910835";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"03fdcb0c";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"1f052408";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"0e001204";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"000908f9";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"ff6608f9";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"003e08f9";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"0307c22c";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"13036514";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"0203bf08";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"0b007804";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"ff8c08f9";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"000d08f9";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"1d027c08";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"0f000604";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"002f08f9";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"00bc08f9";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"000108f9";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"1b025710";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"11006908";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"0c006504";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"006f08f9";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"ff8808f9";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"10004804";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"003108f9";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"00bf08f9";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"1303ff04";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"ff6808f9";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"fff008f9";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"0700f914";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"1cfec804";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"fff908f9";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"00fc1108";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"00fbbc04";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"006408f9";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"ffc108f9";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"01079704";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"00a208f9";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"002908f9";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"0f000808";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"14040004";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"00a908f9";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"ffbf08f9";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"03103e08";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"17f79204";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"007208f9";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"ffaa08f9";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"08003a04";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"ffeb08f9";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"008708f9";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"03fdcb0c";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"1f052408";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"0a003804";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"001109bd";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"ff6709bd";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"003b09bd";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"0307c228";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"13036514";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"0203bf08";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"0e002b04";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"000909bd";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"ff9209bd";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"1d027c08";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"09009b04";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"00bf09bd";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"003a09bd";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"000209bd";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"1b02520c";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"04f92e04";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"ffa409bd";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"04fb1404";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"00a609bd";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"001609bd";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"06fe6f04";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"ff7109bd";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"000009bd";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"0700f914";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"1cfec804";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"fffa09bd";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"07fd7a08";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"08003c04";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"ffc109bd";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"005f09bd";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"01079704";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"009e09bd";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"002e09bd";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"0f00080c";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"0d000904";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"ffd709bd";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"0d00ad04";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"00a909bd";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"003009bd";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"03103e08";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"17f79204";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"006c09bd";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"ffb409bd";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"1e026304";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"ffe809bd";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"008109bd";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"03fca208";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"1f052404";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"ff670a49";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"003c0a49";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"030c2c1c";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"1afa750c";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"19000704";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"ffaa0a49";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"0900e004";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"002b0a49";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"00b60a49";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"1f027b0c";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"00fd1a04";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"ff830a49";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"03033e04";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"ffe10a49";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"003d0a49";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"ff7a0a49";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"19000110";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"1afbf508";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"00fc9e04";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"ffbd0a49";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"00660a49";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"13040004";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"009e0a49";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"00150a49";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"19000308";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"02065904";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"ff7e0a49";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"000f0a49";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"09006104";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"ffe10a49";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"11008004";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"00260a49";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"00840a49";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"03fca208";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"1f052404";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"ff680ad9";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"00350ad9";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"0307c21c";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"0e001d08";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"0003f804";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"ffd10ad9";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"00e50ad9";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"1000560c";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"1af8eb04";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"00690ad9";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"17f73504";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"00150ad9";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"ff910ad9";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"10005804";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"00920ad9";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"fff60ad9";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"1b026a10";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"02045b08";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"0203b504";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"005e0ad9";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"ffa50ad9";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"13040004";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"00970ad9";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"00220ad9";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"17f7e508";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"1b026e04";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"000a0ad9";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"ff5f0ad9";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"03145b08";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"04facb04";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"ffe50ad9";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"00760ad9";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"008a0ad9";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"03fca208";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"1f052404";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"ff690b2d";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"00330b2d";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"03145b1c";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"010e8418";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"1afa7508";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"19000504";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"ffe10b2d";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"008d0b2d";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"19000108";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"12007704";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"004d0b2d";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"ffef0b2d";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"10003d04";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"002f0b2d";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"ff9c0b2d";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"ff920b2d";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"0900eb04";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"008e0b2d";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"00000b2d";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"03fca208";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"1ef9ac04";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"00300bc1";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"ff690bc1";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"030e8430";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"07027d14";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"0e001f08";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"04fca304";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"001c0bc1";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"00b60bc1";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"10004104";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"ff980bc1";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"07ff1604";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"ffab0bc1";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"002e0bc1";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"17f7be0c";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"0f000608";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"0900b504";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"00070bc1";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"ff950bc1";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"00750bc1";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"05f93108";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"08004704";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"ff760bc1";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"ffdf0bc1";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"0d006804";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"00340bc1";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"ffba0bc1";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"10004304";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"008c0bc1";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"0e00330c";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"0c009d04";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"005e0bc1";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"04f92e04";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"000e0bc1";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"ff5e0bc1";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"007b0bc1";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"03fca208";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"0b00b704";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"ff6a0c45";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"00330c45";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"030c2c20";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"0e001d08";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"04fc6804";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"ffce0c45";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"00a10c45";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"0c00b210";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"03003708";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"19000204";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"ff910c45";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"000d0c45";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"04f8fc04";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"ffd00c45";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"00350c45";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"04f94504";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"000b0c45";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"ff7c0c45";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"1900010c";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"020b5c08";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"0b008e04";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"00930c45";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"fff90c45";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"fff10c45";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"19000308";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"1c026b04";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"ff9e0c45";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"ffe60c45";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"0a004804";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"00720c45";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"fff20c45";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"03fca208";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"0b00b704";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"ff6b0cd9";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"002f0cd9";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"030c2c20";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"05f43904";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"ff950cd9";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"05f6980c";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"0208ef08";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"08004204";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"007a0cd9";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"fff80cd9";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"ffa70cd9";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"11023a08";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"03045c04";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"ff910cd9";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"fff80cd9";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"02035004";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"ffe90cd9";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"006c0cd9";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"0900e918";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"0a004d0c";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"05fa8508";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"11006204";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"001c0cd9";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"00910cd9";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"00160cd9";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"03145b08";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"18004504";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"fff10cd9";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"ffba0cd9";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"00560cd9";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"0900eb04";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"ff970cd9";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"0f001104";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"005f0cd9";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"000e0cd9";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"03fdcb0c";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"08002c08";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"1d028404";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"ff9f0d3d";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"00810d3d";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"ff6c0d3d";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"030e8418";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"04f77004";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"ffa90d3d";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"030c2c10";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"11023a08";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"1f025c04";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"00300d3d";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"ffc90d3d";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"1af9e504";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"006f0d3d";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"00070d3d";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"00700d3d";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"10004404";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"007e0d3d";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"16007608";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"04f92e04";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"001e0d3d";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"ff8b0d3d";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"006d0d3d";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"03fca208";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"0f036304";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"ff6d0dc9";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"002a0dc9";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"0307c224";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"0d013b18";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"010c640c";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"17fa7f08";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"0a004504";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"ff760dc9";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"ffe70dc9";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"00190dc9";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"0d002c08";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"12007404";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"007d0dc9";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"ffd70dc9";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"ffa40dc9";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"04fa9604";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"ffc70dc9";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"1d026a04";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"008a0dc9";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"000f0dc9";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"0f000808";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"13040004";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"00870dc9";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"ffd80dc9";
		wait for Clk_period;
		Addr <=  "0001101101001";
		Trees_din <= x"04facb10";
		wait for Clk_period;
		Addr <=  "0001101101010";
		Trees_din <= x"03103e08";
		wait for Clk_period;
		Addr <=  "0001101101011";
		Trees_din <= x"17f79204";
		wait for Clk_period;
		Addr <=  "0001101101100";
		Trees_din <= x"00550dc9";
		wait for Clk_period;
		Addr <=  "0001101101101";
		Trees_din <= x"ffa70dc9";
		wait for Clk_period;
		Addr <=  "0001101101110";
		Trees_din <= x"0900ea04";
		wait for Clk_period;
		Addr <=  "0001101101111";
		Trees_din <= x"005d0dc9";
		wait for Clk_period;
		Addr <=  "0001101110000";
		Trees_din <= x"ffd60dc9";
		wait for Clk_period;
		Addr <=  "0001101110001";
		Trees_din <= x"00690dc9";
		wait for Clk_period;
		Addr <=  "0001101110010";
		Trees_din <= x"03fdcb0c";
		wait for Clk_period;
		Addr <=  "0001101110011";
		Trees_din <= x"08002c08";
		wait for Clk_period;
		Addr <=  "0001101110100";
		Trees_din <= x"1d028404";
		wait for Clk_period;
		Addr <=  "0001101110101";
		Trees_din <= x"ffa80e2d";
		wait for Clk_period;
		Addr <=  "0001101110110";
		Trees_din <= x"00720e2d";
		wait for Clk_period;
		Addr <=  "0001101110111";
		Trees_din <= x"ff6e0e2d";
		wait for Clk_period;
		Addr <=  "0001101111000";
		Trees_din <= x"010e8424";
		wait for Clk_period;
		Addr <=  "0001101111001";
		Trees_din <= x"05ff3b20";
		wait for Clk_period;
		Addr <=  "0001101111010";
		Trees_din <= x"1b026a10";
		wait for Clk_period;
		Addr <=  "0001101111011";
		Trees_din <= x"0307c208";
		wait for Clk_period;
		Addr <=  "0001101111100";
		Trees_din <= x"0f000604";
		wait for Clk_period;
		Addr <=  "0001101111101";
		Trees_din <= x"ffc80e2d";
		wait for Clk_period;
		Addr <=  "0001101111110";
		Trees_din <= x"00570e2d";
		wait for Clk_period;
		Addr <=  "0001101111111";
		Trees_din <= x"14040004";
		wait for Clk_period;
		Addr <=  "0001110000000";
		Trees_din <= x"00780e2d";
		wait for Clk_period;
		Addr <=  "0001110000001";
		Trees_din <= x"fff40e2d";
		wait for Clk_period;
		Addr <=  "0001110000010";
		Trees_din <= x"17f7e908";
		wait for Clk_period;
		Addr <=  "0001110000011";
		Trees_din <= x"04fb6a04";
		wait for Clk_period;
		Addr <=  "0001110000100";
		Trees_din <= x"ff860e2d";
		wait for Clk_period;
		Addr <=  "0001110000101";
		Trees_din <= x"00420e2d";
		wait for Clk_period;
		Addr <=  "0001110000110";
		Trees_din <= x"00fe5f04";
		wait for Clk_period;
		Addr <=  "0001110000111";
		Trees_din <= x"00580e2d";
		wait for Clk_period;
		Addr <=  "0001110001000";
		Trees_din <= x"00060e2d";
		wait for Clk_period;
		Addr <=  "0001110001001";
		Trees_din <= x"ffba0e2d";
		wait for Clk_period;
		Addr <=  "0001110001010";
		Trees_din <= x"ffa20e2d";
		wait for Clk_period;
		Addr <=  "0001110001011";
		Trees_din <= x"03fca208";
		wait for Clk_period;
		Addr <=  "0001110001100";
		Trees_din <= x"1a018704";
		wait for Clk_period;
		Addr <=  "0001110001101";
		Trees_din <= x"ff700ea9";
		wait for Clk_period;
		Addr <=  "0001110001110";
		Trees_din <= x"001f0ea9";
		wait for Clk_period;
		Addr <=  "0001110001111";
		Trees_din <= x"0307c21c";
		wait for Clk_period;
		Addr <=  "0001110010000";
		Trees_din <= x"04f92e04";
		wait for Clk_period;
		Addr <=  "0001110010001";
		Trees_din <= x"ffa30ea9";
		wait for Clk_period;
		Addr <=  "0001110010010";
		Trees_din <= x"1f025208";
		wait for Clk_period;
		Addr <=  "0001110010011";
		Trees_din <= x"06fc5604";
		wait for Clk_period;
		Addr <=  "0001110010100";
		Trees_din <= x"00630ea9";
		wait for Clk_period;
		Addr <=  "0001110010101";
		Trees_din <= x"fff80ea9";
		wait for Clk_period;
		Addr <=  "0001110010110";
		Trees_din <= x"13035c08";
		wait for Clk_period;
		Addr <=  "0001110010111";
		Trees_din <= x"0203bf04";
		wait for Clk_period;
		Addr <=  "0001110011000";
		Trees_din <= x"ffd70ea9";
		wait for Clk_period;
		Addr <=  "0001110011001";
		Trees_din <= x"00470ea9";
		wait for Clk_period;
		Addr <=  "0001110011010";
		Trees_din <= x"0e001704";
		wait for Clk_period;
		Addr <=  "0001110011011";
		Trees_din <= x"002c0ea9";
		wait for Clk_period;
		Addr <=  "0001110011100";
		Trees_din <= x"ff940ea9";
		wait for Clk_period;
		Addr <=  "0001110011101";
		Trees_din <= x"0f000808";
		wait for Clk_period;
		Addr <=  "0001110011110";
		Trees_din <= x"11000404";
		wait for Clk_period;
		Addr <=  "0001110011111";
		Trees_din <= x"ffe50ea9";
		wait for Clk_period;
		Addr <=  "0001110100000";
		Trees_din <= x"007b0ea9";
		wait for Clk_period;
		Addr <=  "0001110100001";
		Trees_din <= x"0f001108";
		wait for Clk_period;
		Addr <=  "0001110100010";
		Trees_din <= x"00fd6604";
		wait for Clk_period;
		Addr <=  "0001110100011";
		Trees_din <= x"ffa70ea9";
		wait for Clk_period;
		Addr <=  "0001110100100";
		Trees_din <= x"00290ea9";
		wait for Clk_period;
		Addr <=  "0001110100101";
		Trees_din <= x"020b5c08";
		wait for Clk_period;
		Addr <=  "0001110100110";
		Trees_din <= x"06faad04";
		wait for Clk_period;
		Addr <=  "0001110100111";
		Trees_din <= x"00730ea9";
		wait for Clk_period;
		Addr <=  "0001110101000";
		Trees_din <= x"00070ea9";
		wait for Clk_period;
		Addr <=  "0001110101001";
		Trees_din <= x"ffb70ea9";
		wait for Clk_period;
		Addr <=  "0001110101010";
		Trees_din <= x"03fca208";
		wait for Clk_period;
		Addr <=  "0001110101011";
		Trees_din <= x"1a018704";
		wait for Clk_period;
		Addr <=  "0001110101100";
		Trees_din <= x"ff720f05";
		wait for Clk_period;
		Addr <=  "0001110101101";
		Trees_din <= x"001c0f05";
		wait for Clk_period;
		Addr <=  "0001110101110";
		Trees_din <= x"010e8424";
		wait for Clk_period;
		Addr <=  "0001110101111";
		Trees_din <= x"0700a210";
		wait for Clk_period;
		Addr <=  "0001110110000";
		Trees_din <= x"06feca0c";
		wait for Clk_period;
		Addr <=  "0001110110001";
		Trees_din <= x"00fc1104";
		wait for Clk_period;
		Addr <=  "0001110110010";
		Trees_din <= x"ffe00f05";
		wait for Clk_period;
		Addr <=  "0001110110011";
		Trees_din <= x"09006104";
		wait for Clk_period;
		Addr <=  "0001110110100";
		Trees_din <= x"ffe60f05";
		wait for Clk_period;
		Addr <=  "0001110110101";
		Trees_din <= x"00670f05";
		wait for Clk_period;
		Addr <=  "0001110110110";
		Trees_din <= x"ffd80f05";
		wait for Clk_period;
		Addr <=  "0001110110111";
		Trees_din <= x"010d2d10";
		wait for Clk_period;
		Addr <=  "0001110111000";
		Trees_din <= x"1303ad08";
		wait for Clk_period;
		Addr <=  "0001110111001";
		Trees_din <= x"0a004b04";
		wait for Clk_period;
		Addr <=  "0001110111010";
		Trees_din <= x"fff80f05";
		wait for Clk_period;
		Addr <=  "0001110111011";
		Trees_din <= x"005b0f05";
		wait for Clk_period;
		Addr <=  "0001110111100";
		Trees_din <= x"16005f04";
		wait for Clk_period;
		Addr <=  "0001110111101";
		Trees_din <= x"00130f05";
		wait for Clk_period;
		Addr <=  "0001110111110";
		Trees_din <= x"ffb70f05";
		wait for Clk_period;
		Addr <=  "0001110111111";
		Trees_din <= x"00530f05";
		wait for Clk_period;
		Addr <=  "0001111000000";
		Trees_din <= x"ffa30f05";
		wait for Clk_period;
		Addr <=  "0001111000001";
		Trees_din <= x"03fdcb08";
		wait for Clk_period;
		Addr <=  "0001111000010";
		Trees_din <= x"08002c04";
		wait for Clk_period;
		Addr <=  "0001111000011";
		Trees_din <= x"000f0f61";
		wait for Clk_period;
		Addr <=  "0001111000100";
		Trees_din <= x"ff730f61";
		wait for Clk_period;
		Addr <=  "0001111000101";
		Trees_din <= x"03145b20";
		wait for Clk_period;
		Addr <=  "0001111000110";
		Trees_din <= x"14021504";
		wait for Clk_period;
		Addr <=  "0001111000111";
		Trees_din <= x"ffb10f61";
		wait for Clk_period;
		Addr <=  "0001111001000";
		Trees_din <= x"1303ad0c";
		wait for Clk_period;
		Addr <=  "0001111001001";
		Trees_din <= x"02020604";
		wait for Clk_period;
		Addr <=  "0001111001010";
		Trees_din <= x"ffac0f61";
		wait for Clk_period;
		Addr <=  "0001111001011";
		Trees_din <= x"09007304";
		wait for Clk_period;
		Addr <=  "0001111001100";
		Trees_din <= x"ffdb0f61";
		wait for Clk_period;
		Addr <=  "0001111001101";
		Trees_din <= x"00510f61";
		wait for Clk_period;
		Addr <=  "0001111001110";
		Trees_din <= x"17f76908";
		wait for Clk_period;
		Addr <=  "0001111001111";
		Trees_din <= x"0d000f04";
		wait for Clk_period;
		Addr <=  "0001111010000";
		Trees_din <= x"ffeb0f61";
		wait for Clk_period;
		Addr <=  "0001111010001";
		Trees_din <= x"00610f61";
		wait for Clk_period;
		Addr <=  "0001111010010";
		Trees_din <= x"15003104";
		wait for Clk_period;
		Addr <=  "0001111010011";
		Trees_din <= x"00250f61";
		wait for Clk_period;
		Addr <=  "0001111010100";
		Trees_din <= x"ffb20f61";
		wait for Clk_period;
		Addr <=  "0001111010101";
		Trees_din <= x"0900eb04";
		wait for Clk_period;
		Addr <=  "0001111010110";
		Trees_din <= x"00740f61";
		wait for Clk_period;
		Addr <=  "0001111010111";
		Trees_din <= x"fff00f61";
		wait for Clk_period;
		Addr <=  "0001111011000";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  4
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"0607fa58";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"0603ba28";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"06034b18";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"0c004608";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"1afc9804";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"00ca0105";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"ff690105";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"1af8f808";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"0b006004";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"00890105";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"ff6f0105";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"1e064004";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"ff570105";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"ffbc0105";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"1af95504";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"00ca0105";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"07ff4304";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"ff5c0105";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"05f88f04";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"00ca0105";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"ff960105";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"0207c514";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"050e2d10";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"0107b308";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"00099604";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"02150105";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"ff840105";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"010dac04";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"00790105";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"ff670105";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"ff660105";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"03f8310c";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"0a005104";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"ff570105";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"000ac704";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"00370105";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"ff9c0105";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"08003e08";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"020be604";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"00f60105";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"ff7e0105";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"0c00bc04";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"ff600105";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"005f0105";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"060e3424";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"020c7118";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"0008520c";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"0504f808";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"010a5104";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"03450105";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"ffa40105";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"00000105";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"000cd308";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"17f75a04";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"01b00105";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"00000105";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"ff8c0105";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"00fe1804";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"015c0105";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"01030104";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"ff680105";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"00370105";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"02116904";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"04530105";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"00370105";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"0606cc58";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"06034b20";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"0c004608";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"1afc3504";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"00d90211";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"ff710211";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"1af8f80c";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"0b006004";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"00880211";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"18016704";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"000d0211";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"ff5f0211";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"06ff0804";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"ff570211";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"03f8f504";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"ff5c0211";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"ff840211";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"0207901c";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"03f7200c";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"1c028608";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"0900e504";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"ff5d0211";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"fff30211";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"00f50211";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"00035a08";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"18001504";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"00950211";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"ff9f0211";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"010bab04";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"01f00211";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"ff810211";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"0b00840c";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"02088c08";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"0b006704";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"00990211";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"ff6e0211";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"ff5a0211";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"0b008708";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"1d026b04";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"01d60211";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"ffa50211";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"08004804";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"ff6b0211";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"00270211";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"020db920";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"0007d414";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"0e001804";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"ff880211";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"050b6008";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"010a5104";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"01a80211";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"fffa0211";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"0b007704";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"ff980211";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"00330211";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"17f73004";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"01530211";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"11021704";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"ff6f0211";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"00ac0211";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"060d0404";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"ff6c0211";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"10004704";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"01610211";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"0c009804";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"00b70211";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"ff8f0211";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"0606cc5c";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"06034b24";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"06fedb0c";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"1af89f08";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"0d001904";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"003e033d";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"ff81033d";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"ff5b033d";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"0c004608";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"17f76c04";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"ffaa033d";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"00ce033d";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"03f8f508";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"1af8f804";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"ffc1033d";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"ff60033d";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"ffde033d";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"ff7a033d";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"0207901c";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"03f7200c";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"0900e304";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"ff61033d";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"0d008504";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"ffc1033d";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"0149033d";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"00035a08";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"18001504";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"007d033d";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"ffa7033d";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"010bab04";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"013c033d";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"ff89033d";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"0b00840c";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"02088c08";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"0900e404";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"ff72033d";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"0096033d";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"ff5f033d";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"0b008708";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"1d026b04";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"016e033d";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"ffab033d";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"08004804";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"ff71033d";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"0026033d";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"020bce18";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"000cd314";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"0900f90c";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"0511b808";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"010ec204";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"0134033d";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"ffaa033d";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"ff9f033d";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"05faad04";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"ff67033d";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"00cc033d";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"ff98033d";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"060d0414";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"0106310c";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"0d015304";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"ff60033d";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"13027e04";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"ffa3033d";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"00cd033d";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"11014804";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"002a033d";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"0127033d";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"0003f80c";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"1303f708";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"07f76704";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"0069033d";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"0154033d";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"fff3033d";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"ffa4033d";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"0606cc4c";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"0603ba24";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"06ffc310";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"1af8f80c";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"15002d04";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"00420449";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"0e003904";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"ff6a0449";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"003c0449";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"ff610449";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"1af8d908";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"14034404";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"ff8b0449";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"01150449";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"0c004604";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"005d0449";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"03f8f504";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"ff680449";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"ff9f0449";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"02076e14";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"03f53404";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"ff720449";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"08004308";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"050e2d04";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"00d30449";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"ff960449";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"03f95e04";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"ff630449";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"00640449";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"03f83104";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"ff640449";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"0b008308";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"11002404";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"009c0449";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"ff6b0449";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"03f92804";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"01360449";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"ffd50449";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"060ba424";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"020c411c";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"12007410";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"15004908";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"1c027804";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"ff7d0449";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"009f0449";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"1101f004";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"01300449";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"00010449";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"11000c04";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"ffac0449";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"04022504";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"01050449";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"ffcd0449";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"18014204";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"ff6d0449";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"00690449";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"02107810";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"15002804";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"fff30449";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"0007c308";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"07f60904";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"004c0449";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"010d0449";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"000d0449";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"06112304";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"ff8f0449";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"00ab0449";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"0604df54";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"06034b2c";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"06fedb0c";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"1af89f08";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"01068104";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"00440575";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"ff910575";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"ff600575";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"03f8e610";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"02010208";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"05f68604";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"00c60575";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"ff8f0575";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"13009f04";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"001e0575";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"ff660575";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"010ac008";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"01089804";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"ff9b0575";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"00590575";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"17fff904";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"ff720575";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"00100575";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"07fedb14";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"17f99808";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"0c00d304";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"ff600575";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"001a0575";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"03f9f508";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"0a004004";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"00380575";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"ff870575";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"00ee0575";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"00035a08";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"17f76804";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"00300575";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"ff750575";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"0900dc08";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"05f56304";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"00c60575";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"ff8a0575";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"01240575";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"0607fa2c";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"0208d41c";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"0202ae0c";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"1403ff04";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"ff750575";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"07008f04";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"00b10575";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"ffa20575";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"08004308";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"000b0d04";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"00fa0575";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"ff900575";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"08004904";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"ff900575";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"00740575";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"0104b104";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"ff630575";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"05f5e004";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"ff7e0575";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"05f6b604";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"010d0575";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"ff9e0575";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"0e001804";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"ff810575";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"0210780c";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"000cd308";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"060ba404";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"008c0575";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"00dd0575";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"ffa10575";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"06112304";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"ff810575";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"00990575";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"0603ba5c";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"06ffc320";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"1af8f80c";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"04ff4b04";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"ff7806e1";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"04006304";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"00c006e1";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"ff9206e1";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"06ff0804";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"ff6206e1";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"0a003c08";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"0a003b04";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"ff8906e1";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"00df06e1";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"0c00f104";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"ff6a06e1";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"003406e1";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"03f8e61c";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"10005610";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"1af95508";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"13028c04";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"00c606e1";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"ff7f06e1";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"08004c04";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"ff6506e1";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"ffd906e1";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"10005808";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"10005704";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"00d906e1";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"003206e1";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"ff7b06e1";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"08003e10";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"010ac008";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"01076204";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"ffb706e1";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"013006e1";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"17f98104";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"ff6f06e1";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"004306e1";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"17fa9408";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"01fc8c04";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"000b06e1";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"ff6206e1";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"0f014604";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"00c306e1";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"ffa406e1";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"06078138";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"03f7de1c";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"0900e310";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"06071308";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"16008f04";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"ff6006e1";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"001106e1";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"0a004a04";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"ff9f06e1";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"00a406e1";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"02073808";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"0e002b04";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"ffa106e1";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"00ef06e1";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"ff7906e1";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"00034410";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"00003a08";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"10004604";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"ff9f06e1";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"00cd06e1";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"0d01d604";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"ff5e06e1";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"007f06e1";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"010bab08";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"00054f04";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"00f106e1";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"003506e1";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"ff8906e1";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"0e001804";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"ff8706e1";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"060ba410";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"1403fe08";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"04022504";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"00a706e1";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"ffd006e1";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"15004804";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"ffb806e1";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"00b906e1";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"16006e08";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"04f8fc04";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"001f06e1";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"00e106e1";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"020a6a04";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"00cd06e1";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"fff106e1";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"0603ba40";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"06fedb0c";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"1af89f08";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"0d003c04";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"00440815";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"ffa10815";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"ff640815";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"03f8e614";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"1af95508";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"0b006704";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"00f30815";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"ff780815";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"13009f04";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"003b0815";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"0c004604";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"00150815";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"ff6e0815";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"08003f10";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"1101d808";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"0a003d04";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"00a70815";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"ff950815";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"0f008104";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"ffe80815";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"01b90815";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"1802e608";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"07036e04";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"ff6d0815";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"00030815";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"19000204";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"ff8f0815";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"00d70815";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"06078134";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"03f7de18";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"0f011d10";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"0c009f08";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"0c008b04";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"ff790815";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"00340815";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"07026504";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"ff660815";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"00080815";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"14034804";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"ffe50815";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"00d20815";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"00034410";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"00003a08";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"1403b704";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"ffa60815";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"00af0815";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"0d01d604";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"ff630815";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"00700815";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"05f40804";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"ff8a0815";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"04035104";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"009d0815";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"ff980815";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"060e3414";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"2003ff04";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"ff650815";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"020db908";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"1403ff04";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"00920815";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"001b0815";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"03f7a104";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"ff8b0815";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"001c0815";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"07f62504";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"00100815";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"0002ed08";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"04f8fc04";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"001a0815";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"00c70815";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"06132b04";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"ffc30815";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"00930815";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"0603ba44";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"06fedb14";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"1af89f08";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"1b027d04";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"ffa80925";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"00410925";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"0209d004";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"ff630925";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"0d01bd04";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"ff790925";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"00380925";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"03f8e61c";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"0201020c";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"05f68604";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"00d20925";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"0900ec04";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"ff7f0925";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"002f0925";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"13028c08";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"13026a04";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"ff860925";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"00b40925";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"04fa2204";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"fff10925";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"ff680925";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"00036a04";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"ff690925";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"010ac008";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"0208ef04";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"00690925";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"ff770925";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"0f00d704";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"ff7b0925";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"00190925";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"060ba424";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"0206d510";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"050e2d0c";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"010dac08";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"03f40604";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"ffae0925";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"00870925";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"ff910925";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"ff880925";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"03f4f104";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"ff650925";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"09005808";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"04010504";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"00fc0925";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"fffc0925";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"0e002f04";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"00270925";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"ffbb0925";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"08004714";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"15002804";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"ffdc0925";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"01faca08";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"0a004804";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"007e0925";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"ff810925";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"07f60904";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"00150925";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"00bd0925";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"00023b04";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"00970925";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"0b007d04";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"ff360925";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"006d0925";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"06031340";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"06fedb14";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"1af89f08";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"0b007204";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"ffad0a31";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"00430a31";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"0209d004";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"ff640a31";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"0d01bd04";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"ff7e0a31";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"003a0a31";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"1100e010";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"02fe5604";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"002f0a31";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"01030108";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"1403fd04";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"00430a31";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"ff870a31";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"ff650a31";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"2004000c";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"03f84004";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"ff7a0a31";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"08004304";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"011c0a31";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"ff8e0a31";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"1af8f808";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"13029b04";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"00db0a31";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"ff920a31";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"08004c04";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"ff850a31";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"00420a31";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"0606cc1c";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"03f5ec08";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"1afa1804";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"ffef0a31";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"ff6f0a31";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"08003304";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"ff750a31";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"08004308";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"10004204";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"ffe10a31";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"006d0a31";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"19002704";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"ff8b0a31";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"007e0a31";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"060e3414";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"2003ff04";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"ff700a31";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"0900f908";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"01ff8f04";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"000b0a31";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"00760a31";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"14040004";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"ff510a31";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"00400a31";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"1101910c";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"00042c08";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"2003fb04";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"00230a31";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"00b70a31";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"00320a31";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"11020108";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"0d00f904";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"00600a31";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"ff730a31";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"008d0a31";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"0602803c";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"06fedb10";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"1af89f04";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"fffa0b35";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"0209d004";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"ff650b35";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"07003204";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"ff820b35";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"00450b35";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"0008d218";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"08003f0c";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"11008f04";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"ff750b35";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"07fe5b04";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"00b60b35";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"ffc90b35";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"01fc8c04";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"00160b35";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"0e004a04";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"ff680b35";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"00220b35";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"1af8f808";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"0b006004";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"00b50b35";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"ff9c0b35";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"0b005104";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"00200b35";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"08004c04";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"ff6d0b35";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"fff10b35";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"06078128";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"03f5ec08";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"1c028704";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"ff6f0b35";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"003a0b35";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"01063110";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"07fe2708";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"0900ea04";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"ff7b0b35";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"00010b35";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"0f000104";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"00970b35";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"ffe50b35";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"010bab08";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"0d000c04";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"ffc20b35";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"00a10b35";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"1f028604";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"ff780b35";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"002e0b35";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"0e001804";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"ff8b0b35";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"02068c0c";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"050b6008";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"00085204";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"00a00b35";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"ffea0b35";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"ffdd0b35";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"0f000f08";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"04ff7404";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"ff9f0b35";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"00510b35";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"2003ff04";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"ffad0b35";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"008c0b35";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"06028034";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"06fedb10";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"1af89f04";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"00010c11";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"0209d004";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"ff660c11";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"0d01bd04";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"ff870c11";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"00480c11";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"20040010";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"1100f304";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"ff730c11";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"03f84004";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"ff860c11";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"1b027a04";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"01180c11";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"ffd40c11";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"0c004604";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"00790c11";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"1af8f808";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"13029b04";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"00ae0c11";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"ff990c11";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"0c00aa04";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"ff670c11";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"ffa40c11";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"060ba424";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"04022518";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"08003108";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"16004804";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"fff10c11";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"ff630c11";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"03f42d08";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"0900d304";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"ff5d0c11";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"ffe20c11";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"2003ff04";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"ff6f0c11";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"003e0c11";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"1dfe9204";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"00950c11";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"21000004";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"ff600c11";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"002a0c11";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"08004710";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"0c00e30c";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"13040008";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"020f5a04";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"009d0c11";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"00230c11";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"00050c11";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"ffcf0c11";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"0001e804";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"00760c11";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"ff970c11";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"06028044";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"06fedb10";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"1af89f04";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"00080cfd";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"0209d004";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"ff670cfd";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"0d01bd04";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"ff8d0cfd";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"00480cfd";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"0008d218";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"08003f0c";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"11008f04";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"ff7d0cfd";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"0700bc04";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"00840cfd";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"ffa80cfd";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"0e004a08";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"01fc8c04";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"002e0cfd";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"ff6c0cfd";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"001e0cfd";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"13029710";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"13026a08";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"0c008804";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"00290cfd";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"ff7c0cfd";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"05f3e104";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"00bf0cfd";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"002b0cfd";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"04054304";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"ff690cfd";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"05f75104";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"ff9d0cfd";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"00410cfd";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"060e341c";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"14013608";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"0f02ac04";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"00de0cfd";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"00150cfd";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"000b6a0c";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"2003ff04";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"ff6a0cfd";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"00034404";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"ffe90cfd";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"00330cfd";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"0d000104";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"002c0cfd";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"ff750cfd";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"1101910c";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"00042c08";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"2003ff04";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"002d0cfd";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"00a40cfd";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"00270cfd";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"11020108";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"05f80604";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"ff960cfd";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"001c0cfd";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"00720cfd";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"06028034";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"06fedb10";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"1af89f04";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"000e0de9";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"0209d004";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"ff680de9";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"0e003a04";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"ff920de9";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"00480de9";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"20040010";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"1100f304";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"ff790de9";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"15003004";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"01240de9";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"04fe1e04";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"00820de9";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"ff7f0de9";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"0c004604";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"00690de9";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"1af8f808";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"13029b04";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"00920de9";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"ffa40de9";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"0c00aa04";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"ff6a0de9";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"ffb30de9";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"060ba424";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"04022518";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"08003108";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"15002a04";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"fff00de9";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"ff6c0de9";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"03f5e508";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"16009604";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"ff980de9";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"008e0de9";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"0c009c04";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"ffe70de9";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"004b0de9";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"1dfe9204";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"00780de9";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"21000004";
		wait for Clk_period;
		Addr <=  "0001101101001";
		Trees_din <= x"ff630de9";
		wait for Clk_period;
		Addr <=  "0001101101010";
		Trees_din <= x"002b0de9";
		wait for Clk_period;
		Addr <=  "0001101101011";
		Trees_din <= x"16006e10";
		wait for Clk_period;
		Addr <=  "0001101101100";
		Trees_din <= x"0c00e30c";
		wait for Clk_period;
		Addr <=  "0001101101101";
		Trees_din <= x"01faca08";
		wait for Clk_period;
		Addr <=  "0001101101110";
		Trees_din <= x"12007904";
		wait for Clk_period;
		Addr <=  "0001101101111";
		Trees_din <= x"007c0de9";
		wait for Clk_period;
		Addr <=  "0001101110000";
		Trees_din <= x"ffea0de9";
		wait for Clk_period;
		Addr <=  "0001101110001";
		Trees_din <= x"00a40de9";
		wait for Clk_period;
		Addr <=  "0001101110010";
		Trees_din <= x"ffcf0de9";
		wait for Clk_period;
		Addr <=  "0001101110011";
		Trees_din <= x"020a6a04";
		wait for Clk_period;
		Addr <=  "0001101110100";
		Trees_din <= x"00880de9";
		wait for Clk_period;
		Addr <=  "0001101110101";
		Trees_din <= x"0001e808";
		wait for Clk_period;
		Addr <=  "0001101110110";
		Trees_din <= x"020f5a04";
		wait for Clk_period;
		Addr <=  "0001101110111";
		Trees_din <= x"00760de9";
		wait for Clk_period;
		Addr <=  "0001101111000";
		Trees_din <= x"ffd80de9";
		wait for Clk_period;
		Addr <=  "0001101111001";
		Trees_din <= x"ff500de9";
		wait for Clk_period;
		Addr <=  "0001101111010";
		Trees_din <= x"06028034";
		wait for Clk_period;
		Addr <=  "0001101111011";
		Trees_din <= x"06fedb10";
		wait for Clk_period;
		Addr <=  "0001101111100";
		Trees_din <= x"1af89f04";
		wait for Clk_period;
		Addr <=  "0001101111101";
		Trees_din <= x"00110eed";
		wait for Clk_period;
		Addr <=  "0001101111110";
		Trees_din <= x"0209d004";
		wait for Clk_period;
		Addr <=  "0001101111111";
		Trees_din <= x"ff690eed";
		wait for Clk_period;
		Addr <=  "0001110000000";
		Trees_din <= x"0e003a04";
		wait for Clk_period;
		Addr <=  "0001110000001";
		Trees_din <= x"ff980eed";
		wait for Clk_period;
		Addr <=  "0001110000010";
		Trees_din <= x"004a0eed";
		wait for Clk_period;
		Addr <=  "0001110000011";
		Trees_din <= x"11008f04";
		wait for Clk_period;
		Addr <=  "0001110000100";
		Trees_din <= x"ff700eed";
		wait for Clk_period;
		Addr <=  "0001110000101";
		Trees_din <= x"08003f10";
		wait for Clk_period;
		Addr <=  "0001110000110";
		Trees_din <= x"00077208";
		wait for Clk_period;
		Addr <=  "0001110000111";
		Trees_din <= x"00062604";
		wait for Clk_period;
		Addr <=  "0001110001000";
		Trees_din <= x"fff50eed";
		wait for Clk_period;
		Addr <=  "0001110001001";
		Trees_din <= x"01120eed";
		wait for Clk_period;
		Addr <=  "0001110001010";
		Trees_din <= x"0b005e04";
		wait for Clk_period;
		Addr <=  "0001110001011";
		Trees_din <= x"00740eed";
		wait for Clk_period;
		Addr <=  "0001110001100";
		Trees_din <= x"ff9d0eed";
		wait for Clk_period;
		Addr <=  "0001110001101";
		Trees_din <= x"0a003c08";
		wait for Clk_period;
		Addr <=  "0001110001110";
		Trees_din <= x"15004004";
		wait for Clk_period;
		Addr <=  "0001110001111";
		Trees_din <= x"ffa70eed";
		wait for Clk_period;
		Addr <=  "0001110010000";
		Trees_din <= x"00970eed";
		wait for Clk_period;
		Addr <=  "0001110010001";
		Trees_din <= x"0f000104";
		wait for Clk_period;
		Addr <=  "0001110010010";
		Trees_din <= x"00270eed";
		wait for Clk_period;
		Addr <=  "0001110010011";
		Trees_din <= x"ff780eed";
		wait for Clk_period;
		Addr <=  "0001110010100";
		Trees_din <= x"06078130";
		wait for Clk_period;
		Addr <=  "0001110010101";
		Trees_din <= x"00034414";
		wait for Clk_period;
		Addr <=  "0001110010110";
		Trees_din <= x"05f6e208";
		wait for Clk_period;
		Addr <=  "0001110010111";
		Trees_din <= x"05f6cc04";
		wait for Clk_period;
		Addr <=  "0001110011000";
		Trees_din <= x"ff9c0eed";
		wait for Clk_period;
		Addr <=  "0001110011001";
		Trees_din <= x"00940eed";
		wait for Clk_period;
		Addr <=  "0001110011010";
		Trees_din <= x"00003a08";
		wait for Clk_period;
		Addr <=  "0001110011011";
		Trees_din <= x"0f000104";
		wait for Clk_period;
		Addr <=  "0001110011100";
		Trees_din <= x"007a0eed";
		wait for Clk_period;
		Addr <=  "0001110011101";
		Trees_din <= x"ffaf0eed";
		wait for Clk_period;
		Addr <=  "0001110011110";
		Trees_din <= x"ff600eed";
		wait for Clk_period;
		Addr <=  "0001110011111";
		Trees_din <= x"03f77e0c";
		wait for Clk_period;
		Addr <=  "0001110100000";
		Trees_din <= x"0f013e08";
		wait for Clk_period;
		Addr <=  "0001110100001";
		Trees_din <= x"00068c04";
		wait for Clk_period;
		Addr <=  "0001110100010";
		Trees_din <= x"ffed0eed";
		wait for Clk_period;
		Addr <=  "0001110100011";
		Trees_din <= x"ff840eed";
		wait for Clk_period;
		Addr <=  "0001110100100";
		Trees_din <= x"008b0eed";
		wait for Clk_period;
		Addr <=  "0001110100101";
		Trees_din <= x"1f026608";
		wait for Clk_period;
		Addr <=  "0001110100110";
		Trees_din <= x"010acf04";
		wait for Clk_period;
		Addr <=  "0001110100111";
		Trees_din <= x"00980eed";
		wait for Clk_period;
		Addr <=  "0001110101000";
		Trees_din <= x"ffa30eed";
		wait for Clk_period;
		Addr <=  "0001110101001";
		Trees_din <= x"19000104";
		wait for Clk_period;
		Addr <=  "0001110101010";
		Trees_din <= x"ff8a0eed";
		wait for Clk_period;
		Addr <=  "0001110101011";
		Trees_din <= x"00240eed";
		wait for Clk_period;
		Addr <=  "0001110101100";
		Trees_din <= x"1404001c";
		wait for Clk_period;
		Addr <=  "0001110101101";
		Trees_din <= x"0f00030c";
		wait for Clk_period;
		Addr <=  "0001110101110";
		Trees_din <= x"0e004508";
		wait for Clk_period;
		Addr <=  "0001110101111";
		Trees_din <= x"060e3404";
		wait for Clk_period;
		Addr <=  "0001110110000";
		Trees_din <= x"ff750eed";
		wait for Clk_period;
		Addr <=  "0001110110001";
		Trees_din <= x"00570eed";
		wait for Clk_period;
		Addr <=  "0001110110010";
		Trees_din <= x"007a0eed";
		wait for Clk_period;
		Addr <=  "0001110110011";
		Trees_din <= x"04fe1308";
		wait for Clk_period;
		Addr <=  "0001110110100";
		Trees_din <= x"15003504";
		wait for Clk_period;
		Addr <=  "0001110110101";
		Trees_din <= x"fff60eed";
		wait for Clk_period;
		Addr <=  "0001110110110";
		Trees_din <= x"009b0eed";
		wait for Clk_period;
		Addr <=  "0001110110111";
		Trees_din <= x"07fd9204";
		wait for Clk_period;
		Addr <=  "0001110111000";
		Trees_din <= x"004b0eed";
		wait for Clk_period;
		Addr <=  "0001110111001";
		Trees_din <= x"ffae0eed";
		wait for Clk_period;
		Addr <=  "0001110111010";
		Trees_din <= x"00ae0eed";
		wait for Clk_period;
		Addr <=  "0001110111011";
		Trees_din <= x"06013328";
		wait for Clk_period;
		Addr <=  "0001110111100";
		Trees_din <= x"05f5bf10";
		wait for Clk_period;
		Addr <=  "0001110111101";
		Trees_din <= x"0200ea04";
		wait for Clk_period;
		Addr <=  "0001110111110";
		Trees_din <= x"00170fd1";
		wait for Clk_period;
		Addr <=  "0001110111111";
		Trees_din <= x"00058708";
		wait for Clk_period;
		Addr <=  "0001111000000";
		Trees_din <= x"03f98c04";
		wait for Clk_period;
		Addr <=  "0001111000001";
		Trees_din <= x"00470fd1";
		wait for Clk_period;
		Addr <=  "0001111000010";
		Trees_din <= x"ff830fd1";
		wait for Clk_period;
		Addr <=  "0001111000011";
		Trees_din <= x"ff690fd1";
		wait for Clk_period;
		Addr <=  "0001111000100";
		Trees_din <= x"1100e004";
		wait for Clk_period;
		Addr <=  "0001111000101";
		Trees_din <= x"ff700fd1";
		wait for Clk_period;
		Addr <=  "0001111000110";
		Trees_din <= x"04fc7e04";
		wait for Clk_period;
		Addr <=  "0001111000111";
		Trees_din <= x"ff760fd1";
		wait for Clk_period;
		Addr <=  "0001111001000";
		Trees_din <= x"04ff9108";
		wait for Clk_period;
		Addr <=  "0001111001001";
		Trees_din <= x"02044d04";
		wait for Clk_period;
		Addr <=  "0001111001010";
		Trees_din <= x"ff920fd1";
		wait for Clk_period;
		Addr <=  "0001111001011";
		Trees_din <= x"00d60fd1";
		wait for Clk_period;
		Addr <=  "0001111001100";
		Trees_din <= x"18003604";
		wait for Clk_period;
		Addr <=  "0001111001101";
		Trees_din <= x"00380fd1";
		wait for Clk_period;
		Addr <=  "0001111001110";
		Trees_din <= x"ff790fd1";
		wait for Clk_period;
		Addr <=  "0001111001111";
		Trees_din <= x"14013610";
		wait for Clk_period;
		Addr <=  "0001111010000";
		Trees_din <= x"1101d008";
		wait for Clk_period;
		Addr <=  "0001111010001";
		Trees_din <= x"1303e004";
		wait for Clk_period;
		Addr <=  "0001111010010";
		Trees_din <= x"ffe70fd1";
		wait for Clk_period;
		Addr <=  "0001111010011";
		Trees_din <= x"004d0fd1";
		wait for Clk_period;
		Addr <=  "0001111010100";
		Trees_din <= x"0207ba04";
		wait for Clk_period;
		Addr <=  "0001111010101";
		Trees_din <= x"00470fd1";
		wait for Clk_period;
		Addr <=  "0001111010110";
		Trees_din <= x"01150fd1";
		wait for Clk_period;
		Addr <=  "0001111010111";
		Trees_din <= x"0606cc1c";
		wait for Clk_period;
		Addr <=  "0001111011000";
		Trees_din <= x"0900d510";
		wait for Clk_period;
		Addr <=  "0001111011001";
		Trees_din <= x"07f73f08";
		wait for Clk_period;
		Addr <=  "0001111011010";
		Trees_din <= x"09009104";
		wait for Clk_period;
		Addr <=  "0001111011011";
		Trees_din <= x"00bd0fd1";
		wait for Clk_period;
		Addr <=  "0001111011100";
		Trees_din <= x"000b0fd1";
		wait for Clk_period;
		Addr <=  "0001111011101";
		Trees_din <= x"17f71104";
		wait for Clk_period;
		Addr <=  "0001111011110";
		Trees_din <= x"00150fd1";
		wait for Clk_period;
		Addr <=  "0001111011111";
		Trees_din <= x"ff940fd1";
		wait for Clk_period;
		Addr <=  "0001111100000";
		Trees_din <= x"05f4c904";
		wait for Clk_period;
		Addr <=  "0001111100001";
		Trees_din <= x"ff800fd1";
		wait for Clk_period;
		Addr <=  "0001111100010";
		Trees_din <= x"0003f804";
		wait for Clk_period;
		Addr <=  "0001111100011";
		Trees_din <= x"ffce0fd1";
		wait for Clk_period;
		Addr <=  "0001111100100";
		Trees_din <= x"00580fd1";
		wait for Clk_period;
		Addr <=  "0001111100101";
		Trees_din <= x"0106d810";
		wait for Clk_period;
		Addr <=  "0001111100110";
		Trees_din <= x"060a0b08";
		wait for Clk_period;
		Addr <=  "0001111100111";
		Trees_din <= x"0d000c04";
		wait for Clk_period;
		Addr <=  "0001111101000";
		Trees_din <= x"00710fd1";
		wait for Clk_period;
		Addr <=  "0001111101001";
		Trees_din <= x"ffbf0fd1";
		wait for Clk_period;
		Addr <=  "0001111101010";
		Trees_din <= x"020a8004";
		wait for Clk_period;
		Addr <=  "0001111101011";
		Trees_din <= x"007a0fd1";
		wait for Clk_period;
		Addr <=  "0001111101100";
		Trees_din <= x"00040fd1";
		wait for Clk_period;
		Addr <=  "0001111101101";
		Trees_din <= x"12007408";
		wait for Clk_period;
		Addr <=  "0001111101110";
		Trees_din <= x"0a004604";
		wait for Clk_period;
		Addr <=  "0001111101111";
		Trees_din <= x"ff680fd1";
		wait for Clk_period;
		Addr <=  "0001111110000";
		Trees_din <= x"00810fd1";
		wait for Clk_period;
		Addr <=  "0001111110001";
		Trees_din <= x"0c00dd04";
		wait for Clk_period;
		Addr <=  "0001111110010";
		Trees_din <= x"00cd0fd1";
		wait for Clk_period;
		Addr <=  "0001111110011";
		Trees_din <= x"fff50fd1";
		wait for Clk_period;
		Addr <=  "0001111110100";
		Trees_din <= x"0601332c";
		wait for Clk_period;
		Addr <=  "0001111110101";
		Trees_din <= x"05f5bf10";
		wait for Clk_period;
		Addr <=  "0001111110110";
		Trees_din <= x"0200ea04";
		wait for Clk_period;
		Addr <=  "0001111110111";
		Trees_din <= x"001910ad";
		wait for Clk_period;
		Addr <=  "0001111111000";
		Trees_din <= x"00058708";
		wait for Clk_period;
		Addr <=  "0001111111001";
		Trees_din <= x"05f3b604";
		wait for Clk_period;
		Addr <=  "0001111111010";
		Trees_din <= x"004510ad";
		wait for Clk_period;
		Addr <=  "0001111111011";
		Trees_din <= x"ff8710ad";
		wait for Clk_period;
		Addr <=  "0001111111100";
		Trees_din <= x"ff6b10ad";
		wait for Clk_period;
		Addr <=  "0001111111101";
		Trees_din <= x"05f7a710";
		wait for Clk_period;
		Addr <=  "0001111111110";
		Trees_din <= x"1100e004";
		wait for Clk_period;
		Addr <=  "0001111111111";
		Trees_din <= x"ff7e10ad";
		wait for Clk_period;
		Addr <=  "0010000000000";
		Trees_din <= x"03f84a04";
		wait for Clk_period;
		Addr <=  "0010000000001";
		Trees_din <= x"ff9110ad";
		wait for Clk_period;
		Addr <=  "0010000000010";
		Trees_din <= x"04fc7e04";
		wait for Clk_period;
		Addr <=  "0010000000011";
		Trees_din <= x"ff9810ad";
		wait for Clk_period;
		Addr <=  "0010000000100";
		Trees_din <= x"009810ad";
		wait for Clk_period;
		Addr <=  "0010000000101";
		Trees_din <= x"0c00f108";
		wait for Clk_period;
		Addr <=  "0010000000110";
		Trees_din <= x"11030804";
		wait for Clk_period;
		Addr <=  "0010000000111";
		Trees_din <= x"ff6e10ad";
		wait for Clk_period;
		Addr <=  "0010000001000";
		Trees_din <= x"ffff10ad";
		wait for Clk_period;
		Addr <=  "0010000001001";
		Trees_din <= x"003910ad";
		wait for Clk_period;
		Addr <=  "0010000001010";
		Trees_din <= x"1401360c";
		wait for Clk_period;
		Addr <=  "0010000001011";
		Trees_din <= x"03f86708";
		wait for Clk_period;
		Addr <=  "0010000001100";
		Trees_din <= x"00055e04";
		wait for Clk_period;
		Addr <=  "0010000001101";
		Trees_din <= x"004110ad";
		wait for Clk_period;
		Addr <=  "0010000001110";
		Trees_din <= x"ffeb10ad";
		wait for Clk_period;
		Addr <=  "0010000001111";
		Trees_din <= x"00d510ad";
		wait for Clk_period;
		Addr <=  "0010000010000";
		Trees_din <= x"0606cc1c";
		wait for Clk_period;
		Addr <=  "0010000010001";
		Trees_din <= x"0e003910";
		wait for Clk_period;
		Addr <=  "0010000010010";
		Trees_din <= x"16006008";
		wait for Clk_period;
		Addr <=  "0010000010011";
		Trees_din <= x"05f6d304";
		wait for Clk_period;
		Addr <=  "0010000010100";
		Trees_din <= x"ffd510ad";
		wait for Clk_period;
		Addr <=  "0010000010101";
		Trees_din <= x"ff6e10ad";
		wait for Clk_period;
		Addr <=  "0010000010110";
		Trees_din <= x"0003f804";
		wait for Clk_period;
		Addr <=  "0010000010111";
		Trees_din <= x"ffbf10ad";
		wait for Clk_period;
		Addr <=  "0010000011000";
		Trees_din <= x"005310ad";
		wait for Clk_period;
		Addr <=  "0010000011001";
		Trees_din <= x"02035008";
		wait for Clk_period;
		Addr <=  "0010000011010";
		Trees_din <= x"0a004404";
		wait for Clk_period;
		Addr <=  "0010000011011";
		Trees_din <= x"005010ad";
		wait for Clk_period;
		Addr <=  "0010000011100";
		Trees_din <= x"ffd710ad";
		wait for Clk_period;
		Addr <=  "0010000011101";
		Trees_din <= x"ff6610ad";
		wait for Clk_period;
		Addr <=  "0010000011110";
		Trees_din <= x"00ff630c";
		wait for Clk_period;
		Addr <=  "0010000011111";
		Trees_din <= x"05075f08";
		wait for Clk_period;
		Addr <=  "0010000100000";
		Trees_din <= x"0400f704";
		wait for Clk_period;
		Addr <=  "0010000100001";
		Trees_din <= x"009710ad";
		wait for Clk_period;
		Addr <=  "0010000100010";
		Trees_din <= x"001810ad";
		wait for Clk_period;
		Addr <=  "0010000100011";
		Trees_din <= x"ffce10ad";
		wait for Clk_period;
		Addr <=  "0010000100100";
		Trees_din <= x"0106d808";
		wait for Clk_period;
		Addr <=  "0010000100101";
		Trees_din <= x"02068c04";
		wait for Clk_period;
		Addr <=  "0010000100110";
		Trees_din <= x"005910ad";
		wait for Clk_period;
		Addr <=  "0010000100111";
		Trees_din <= x"ffdc10ad";
		wait for Clk_period;
		Addr <=  "0010000101000";
		Trees_din <= x"12007404";
		wait for Clk_period;
		Addr <=  "0010000101001";
		Trees_din <= x"ffc810ad";
		wait for Clk_period;
		Addr <=  "0010000101010";
		Trees_din <= x"00a510ad";
		wait for Clk_period;
		Addr <=  "0010000101011";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0010000101100";
		Trees_din <= x"0601332c";
		wait for Clk_period;
		Addr <=  "0010000101101";
		Trees_din <= x"1100e004";
		wait for Clk_period;
		Addr <=  "0010000101110";
		Trees_din <= x"ff6d118d";
		wait for Clk_period;
		Addr <=  "0010000101111";
		Trees_din <= x"08003f1c";
		wait for Clk_period;
		Addr <=  "0010000110000";
		Trees_din <= x"0b006e10";
		wait for Clk_period;
		Addr <=  "0010000110001";
		Trees_din <= x"0b006d08";
		wait for Clk_period;
		Addr <=  "0010000110010";
		Trees_din <= x"0b006504";
		wait for Clk_period;
		Addr <=  "0010000110011";
		Trees_din <= x"0091118d";
		wait for Clk_period;
		Addr <=  "0010000110100";
		Trees_din <= x"ff8e118d";
		wait for Clk_period;
		Addr <=  "0010000110101";
		Trees_din <= x"0d00d604";
		wait for Clk_period;
		Addr <=  "0010000110110";
		Trees_din <= x"005d118d";
		wait for Clk_period;
		Addr <=  "0010000110111";
		Trees_din <= x"015d118d";
		wait for Clk_period;
		Addr <=  "0010000111000";
		Trees_din <= x"0c00d304";
		wait for Clk_period;
		Addr <=  "0010000111001";
		Trees_din <= x"ff73118d";
		wait for Clk_period;
		Addr <=  "0010000111010";
		Trees_din <= x"0108e504";
		wait for Clk_period;
		Addr <=  "0010000111011";
		Trees_din <= x"00cc118d";
		wait for Clk_period;
		Addr <=  "0010000111100";
		Trees_din <= x"ffc4118d";
		wait for Clk_period;
		Addr <=  "0010000111101";
		Trees_din <= x"03028708";
		wait for Clk_period;
		Addr <=  "0010000111110";
		Trees_din <= x"0e004a04";
		wait for Clk_period;
		Addr <=  "0010000111111";
		Trees_din <= x"ff6d118d";
		wait for Clk_period;
		Addr <=  "0010001000000";
		Trees_din <= x"000b118d";
		wait for Clk_period;
		Addr <=  "0010001000001";
		Trees_din <= x"001d118d";
		wait for Clk_period;
		Addr <=  "0010001000010";
		Trees_din <= x"1401360c";
		wait for Clk_period;
		Addr <=  "0010001000011";
		Trees_din <= x"04ffc904";
		wait for Clk_period;
		Addr <=  "0010001000100";
		Trees_din <= x"fffd118d";
		wait for Clk_period;
		Addr <=  "0010001000101";
		Trees_din <= x"1101d004";
		wait for Clk_period;
		Addr <=  "0010001000110";
		Trees_din <= x"001b118d";
		wait for Clk_period;
		Addr <=  "0010001000111";
		Trees_din <= x"00de118d";
		wait for Clk_period;
		Addr <=  "0010001001000";
		Trees_din <= x"0604df20";
		wait for Clk_period;
		Addr <=  "0010001001001";
		Trees_din <= x"07fedb10";
		wait for Clk_period;
		Addr <=  "0010001001010";
		Trees_din <= x"13028c08";
		wait for Clk_period;
		Addr <=  "0010001001011";
		Trees_din <= x"13026a04";
		wait for Clk_period;
		Addr <=  "0010001001100";
		Trees_din <= x"ffa1118d";
		wait for Clk_period;
		Addr <=  "0010001001101";
		Trees_din <= x"00d8118d";
		wait for Clk_period;
		Addr <=  "0010001001110";
		Trees_din <= x"03fab204";
		wait for Clk_period;
		Addr <=  "0010001001111";
		Trees_din <= x"ff76118d";
		wait for Clk_period;
		Addr <=  "0010001010000";
		Trees_din <= x"0018118d";
		wait for Clk_period;
		Addr <=  "0010001010001";
		Trees_din <= x"0700e908";
		wait for Clk_period;
		Addr <=  "0010001010010";
		Trees_din <= x"13035c04";
		wait for Clk_period;
		Addr <=  "0010001010011";
		Trees_din <= x"ff9b118d";
		wait for Clk_period;
		Addr <=  "0010001010100";
		Trees_din <= x"00b4118d";
		wait for Clk_period;
		Addr <=  "0010001010101";
		Trees_din <= x"0b006f04";
		wait for Clk_period;
		Addr <=  "0010001010110";
		Trees_din <= x"000f118d";
		wait for Clk_period;
		Addr <=  "0010001010111";
		Trees_din <= x"ff85118d";
		wait for Clk_period;
		Addr <=  "0010001011000";
		Trees_din <= x"00fe1808";
		wait for Clk_period;
		Addr <=  "0010001011001";
		Trees_din <= x"06099f04";
		wait for Clk_period;
		Addr <=  "0010001011010";
		Trees_din <= x"000c118d";
		wait for Clk_period;
		Addr <=  "0010001011011";
		Trees_din <= x"008b118d";
		wait for Clk_period;
		Addr <=  "0010001011100";
		Trees_din <= x"05f6ed08";
		wait for Clk_period;
		Addr <=  "0010001011101";
		Trees_din <= x"0106d804";
		wait for Clk_period;
		Addr <=  "0010001011110";
		Trees_din <= x"0000118d";
		wait for Clk_period;
		Addr <=  "0010001011111";
		Trees_din <= x"0088118d";
		wait for Clk_period;
		Addr <=  "0010001100000";
		Trees_din <= x"15004804";
		wait for Clk_period;
		Addr <=  "0010001100001";
		Trees_din <= x"ffdc118d";
		wait for Clk_period;
		Addr <=  "0010001100010";
		Trees_din <= x"0062118d";
		wait for Clk_period;
		Addr <=  "0010001100011";
		Trees_din <= x"06013328";
		wait for Clk_period;
		Addr <=  "0010001100100";
		Trees_din <= x"1100e004";
		wait for Clk_period;
		Addr <=  "0010001100101";
		Trees_din <= x"ff6e1261";
		wait for Clk_period;
		Addr <=  "0010001100110";
		Trees_din <= x"08003f18";
		wait for Clk_period;
		Addr <=  "0010001100111";
		Trees_din <= x"0b006e0c";
		wait for Clk_period;
		Addr <=  "0010001101000";
		Trees_din <= x"06fedb04";
		wait for Clk_period;
		Addr <=  "0010001101001";
		Trees_din <= x"ffa21261";
		wait for Clk_period;
		Addr <=  "0010001101010";
		Trees_din <= x"00076404";
		wait for Clk_period;
		Addr <=  "0010001101011";
		Trees_din <= x"00f01261";
		wait for Clk_period;
		Addr <=  "0010001101100";
		Trees_din <= x"000c1261";
		wait for Clk_period;
		Addr <=  "0010001101101";
		Trees_din <= x"0c00d304";
		wait for Clk_period;
		Addr <=  "0010001101110";
		Trees_din <= x"ff761261";
		wait for Clk_period;
		Addr <=  "0010001101111";
		Trees_din <= x"0d00e904";
		wait for Clk_period;
		Addr <=  "0010001110000";
		Trees_din <= x"009d1261";
		wait for Clk_period;
		Addr <=  "0010001110001";
		Trees_din <= x"ff9f1261";
		wait for Clk_period;
		Addr <=  "0010001110010";
		Trees_din <= x"03028708";
		wait for Clk_period;
		Addr <=  "0010001110011";
		Trees_din <= x"0e004a04";
		wait for Clk_period;
		Addr <=  "0010001110100";
		Trees_din <= x"ff6e1261";
		wait for Clk_period;
		Addr <=  "0010001110101";
		Trees_din <= x"000c1261";
		wait for Clk_period;
		Addr <=  "0010001110110";
		Trees_din <= x"001d1261";
		wait for Clk_period;
		Addr <=  "0010001110111";
		Trees_din <= x"1401360c";
		wait for Clk_period;
		Addr <=  "0010001111000";
		Trees_din <= x"04ffc904";
		wait for Clk_period;
		Addr <=  "0010001111001";
		Trees_din <= x"fffa1261";
		wait for Clk_period;
		Addr <=  "0010001111010";
		Trees_din <= x"03f86704";
		wait for Clk_period;
		Addr <=  "0010001111011";
		Trees_din <= x"00261261";
		wait for Clk_period;
		Addr <=  "0010001111100";
		Trees_din <= x"00c81261";
		wait for Clk_period;
		Addr <=  "0010001111101";
		Trees_din <= x"060ba41c";
		wait for Clk_period;
		Addr <=  "0010001111110";
		Trees_din <= x"0207c50c";
		wait for Clk_period;
		Addr <=  "0010001111111";
		Trees_din <= x"0401c208";
		wait for Clk_period;
		Addr <=  "0010010000000";
		Trees_din <= x"04ffe504";
		wait for Clk_period;
		Addr <=  "0010010000001";
		Trees_din <= x"000b1261";
		wait for Clk_period;
		Addr <=  "0010010000010";
		Trees_din <= x"00871261";
		wait for Clk_period;
		Addr <=  "0010010000011";
		Trees_din <= x"ff711261";
		wait for Clk_period;
		Addr <=  "0010010000100";
		Trees_din <= x"09005808";
		wait for Clk_period;
		Addr <=  "0010010000101";
		Trees_din <= x"01041e04";
		wait for Clk_period;
		Addr <=  "0010010000110";
		Trees_din <= x"00901261";
		wait for Clk_period;
		Addr <=  "0010010000111";
		Trees_din <= x"fffd1261";
		wait for Clk_period;
		Addr <=  "0010010001000";
		Trees_din <= x"0106d804";
		wait for Clk_period;
		Addr <=  "0010010001001";
		Trees_din <= x"ffab1261";
		wait for Clk_period;
		Addr <=  "0010010001010";
		Trees_din <= x"00041261";
		wait for Clk_period;
		Addr <=  "0010010001011";
		Trees_din <= x"16006e0c";
		wait for Clk_period;
		Addr <=  "0010010001100";
		Trees_din <= x"04fa3304";
		wait for Clk_period;
		Addr <=  "0010010001101";
		Trees_din <= x"ffe51261";
		wait for Clk_period;
		Addr <=  "0010010001110";
		Trees_din <= x"08003704";
		wait for Clk_period;
		Addr <=  "0010010001111";
		Trees_din <= x"00271261";
		wait for Clk_period;
		Addr <=  "0010010010000";
		Trees_din <= x"00931261";
		wait for Clk_period;
		Addr <=  "0010010010001";
		Trees_din <= x"16007908";
		wait for Clk_period;
		Addr <=  "0010010010010";
		Trees_din <= x"0e003804";
		wait for Clk_period;
		Addr <=  "0010010010011";
		Trees_din <= x"ff7e1261";
		wait for Clk_period;
		Addr <=  "0010010010100";
		Trees_din <= x"00021261";
		wait for Clk_period;
		Addr <=  "0010010010101";
		Trees_din <= x"17f7e704";
		wait for Clk_period;
		Addr <=  "0010010010110";
		Trees_din <= x"00691261";
		wait for Clk_period;
		Addr <=  "0010010010111";
		Trees_din <= x"001f1261";
		wait for Clk_period;
		Addr <=  "0010010011000";
		Trees_din <= x"06fedb0c";
		wait for Clk_period;
		Addr <=  "0010010011001";
		Trees_din <= x"01068108";
		wait for Clk_period;
		Addr <=  "0010010011010";
		Trees_din <= x"05f6ed04";
		wait for Clk_period;
		Addr <=  "0010010011011";
		Trees_din <= x"006f12fd";
		wait for Clk_period;
		Addr <=  "0010010011100";
		Trees_din <= x"ff8f12fd";
		wait for Clk_period;
		Addr <=  "0010010011101";
		Trees_din <= x"ff6f12fd";
		wait for Clk_period;
		Addr <=  "0010010011110";
		Trees_din <= x"00099624";
		wait for Clk_period;
		Addr <=  "0010010011111";
		Trees_din <= x"010e7620";
		wait for Clk_period;
		Addr <=  "0010010100000";
		Trees_din <= x"0700e910";
		wait for Clk_period;
		Addr <=  "0010010100001";
		Trees_din <= x"02068c08";
		wait for Clk_period;
		Addr <=  "0010010100010";
		Trees_din <= x"05f75104";
		wait for Clk_period;
		Addr <=  "0010010100011";
		Trees_din <= x"00cf12fd";
		wait for Clk_period;
		Addr <=  "0010010100100";
		Trees_din <= x"002112fd";
		wait for Clk_period;
		Addr <=  "0010010100101";
		Trees_din <= x"00094404";
		wait for Clk_period;
		Addr <=  "0010010100110";
		Trees_din <= x"000312fd";
		wait for Clk_period;
		Addr <=  "0010010100111";
		Trees_din <= x"009b12fd";
		wait for Clk_period;
		Addr <=  "0010010101000";
		Trees_din <= x"06058308";
		wait for Clk_period;
		Addr <=  "0010010101001";
		Trees_din <= x"01fe5404";
		wait for Clk_period;
		Addr <=  "0010010101010";
		Trees_din <= x"003c12fd";
		wait for Clk_period;
		Addr <=  "0010010101011";
		Trees_din <= x"ff8412fd";
		wait for Clk_period;
		Addr <=  "0010010101100";
		Trees_din <= x"04fe0304";
		wait for Clk_period;
		Addr <=  "0010010101101";
		Trees_din <= x"006212fd";
		wait for Clk_period;
		Addr <=  "0010010101110";
		Trees_din <= x"ffa712fd";
		wait for Clk_period;
		Addr <=  "0010010101111";
		Trees_din <= x"ff8012fd";
		wait for Clk_period;
		Addr <=  "0010010110000";
		Trees_din <= x"1302970c";
		wait for Clk_period;
		Addr <=  "0010010110001";
		Trees_din <= x"13026a08";
		wait for Clk_period;
		Addr <=  "0010010110010";
		Trees_din <= x"1c025a04";
		wait for Clk_period;
		Addr <=  "0010010110011";
		Trees_din <= x"006512fd";
		wait for Clk_period;
		Addr <=  "0010010110100";
		Trees_din <= x"ff8c12fd";
		wait for Clk_period;
		Addr <=  "0010010110101";
		Trees_din <= x"00ae12fd";
		wait for Clk_period;
		Addr <=  "0010010110110";
		Trees_din <= x"0a003e0c";
		wait for Clk_period;
		Addr <=  "0010010110111";
		Trees_din <= x"0403e708";
		wait for Clk_period;
		Addr <=  "0010010111000";
		Trees_din <= x"18015104";
		wait for Clk_period;
		Addr <=  "0010010111001";
		Trees_din <= x"ff9812fd";
		wait for Clk_period;
		Addr <=  "0010010111010";
		Trees_din <= x"fffe12fd";
		wait for Clk_period;
		Addr <=  "0010010111011";
		Trees_din <= x"006012fd";
		wait for Clk_period;
		Addr <=  "0010010111100";
		Trees_din <= x"05f19304";
		wait for Clk_period;
		Addr <=  "0010010111101";
		Trees_din <= x"fffe12fd";
		wait for Clk_period;
		Addr <=  "0010010111110";
		Trees_din <= x"ff6b12fd";
		wait for Clk_period;
		Addr <=  "0010010111111";
		Trees_din <= x"06013328";
		wait for Clk_period;
		Addr <=  "0010011000000";
		Trees_din <= x"1100e004";
		wait for Clk_period;
		Addr <=  "0010011000001";
		Trees_din <= x"ff7113c9";
		wait for Clk_period;
		Addr <=  "0010011000010";
		Trees_din <= x"08003f18";
		wait for Clk_period;
		Addr <=  "0010011000011";
		Trees_din <= x"0b006e0c";
		wait for Clk_period;
		Addr <=  "0010011000100";
		Trees_din <= x"0b006d08";
		wait for Clk_period;
		Addr <=  "0010011000101";
		Trees_din <= x"12006f04";
		wait for Clk_period;
		Addr <=  "0010011000110";
		Trees_din <= x"007313c9";
		wait for Clk_period;
		Addr <=  "0010011000111";
		Trees_din <= x"ff9413c9";
		wait for Clk_period;
		Addr <=  "0010011001000";
		Trees_din <= x"00d513c9";
		wait for Clk_period;
		Addr <=  "0010011001001";
		Trees_din <= x"15003008";
		wait for Clk_period;
		Addr <=  "0010011001010";
		Trees_din <= x"15002c04";
		wait for Clk_period;
		Addr <=  "0010011001011";
		Trees_din <= x"ffc113c9";
		wait for Clk_period;
		Addr <=  "0010011001100";
		Trees_din <= x"00a513c9";
		wait for Clk_period;
		Addr <=  "0010011001101";
		Trees_din <= x"ff7a13c9";
		wait for Clk_period;
		Addr <=  "0010011001110";
		Trees_din <= x"03028708";
		wait for Clk_period;
		Addr <=  "0010011001111";
		Trees_din <= x"0d037604";
		wait for Clk_period;
		Addr <=  "0010011010000";
		Trees_din <= x"ff7213c9";
		wait for Clk_period;
		Addr <=  "0010011010001";
		Trees_din <= x"001013c9";
		wait for Clk_period;
		Addr <=  "0010011010010";
		Trees_din <= x"002613c9";
		wait for Clk_period;
		Addr <=  "0010011010011";
		Trees_din <= x"2003ff08";
		wait for Clk_period;
		Addr <=  "0010011010100";
		Trees_din <= x"03f66c04";
		wait for Clk_period;
		Addr <=  "0010011010101";
		Trees_din <= x"ffea13c9";
		wait for Clk_period;
		Addr <=  "0010011010110";
		Trees_din <= x"ff8413c9";
		wait for Clk_period;
		Addr <=  "0010011010111";
		Trees_din <= x"20040018";
		wait for Clk_period;
		Addr <=  "0010011011000";
		Trees_din <= x"0e003810";
		wait for Clk_period;
		Addr <=  "0010011011001";
		Trees_din <= x"0a004108";
		wait for Clk_period;
		Addr <=  "0010011011010";
		Trees_din <= x"06078104";
		wait for Clk_period;
		Addr <=  "0010011011011";
		Trees_din <= x"ff9913c9";
		wait for Clk_period;
		Addr <=  "0010011011100";
		Trees_din <= x"006b13c9";
		wait for Clk_period;
		Addr <=  "0010011011101";
		Trees_din <= x"0a005204";
		wait for Clk_period;
		Addr <=  "0010011011110";
		Trees_din <= x"009813c9";
		wait for Clk_period;
		Addr <=  "0010011011111";
		Trees_din <= x"ffe813c9";
		wait for Clk_period;
		Addr <=  "0010011100000";
		Trees_din <= x"0206ab04";
		wait for Clk_period;
		Addr <=  "0010011100001";
		Trees_din <= x"002913c9";
		wait for Clk_period;
		Addr <=  "0010011100010";
		Trees_din <= x"ff9313c9";
		wait for Clk_period;
		Addr <=  "0010011100011";
		Trees_din <= x"0b007a10";
		wait for Clk_period;
		Addr <=  "0010011100100";
		Trees_din <= x"12007908";
		wait for Clk_period;
		Addr <=  "0010011100101";
		Trees_din <= x"060ab504";
		wait for Clk_period;
		Addr <=  "0010011100110";
		Trees_din <= x"ffe913c9";
		wait for Clk_period;
		Addr <=  "0010011100111";
		Trees_din <= x"005f13c9";
		wait for Clk_period;
		Addr <=  "0010011101000";
		Trees_din <= x"03f64204";
		wait for Clk_period;
		Addr <=  "0010011101001";
		Trees_din <= x"ffba13c9";
		wait for Clk_period;
		Addr <=  "0010011101010";
		Trees_din <= x"008e13c9";
		wait for Clk_period;
		Addr <=  "0010011101011";
		Trees_din <= x"16006e08";
		wait for Clk_period;
		Addr <=  "0010011101100";
		Trees_din <= x"0a004104";
		wait for Clk_period;
		Addr <=  "0010011101101";
		Trees_din <= x"ff8c13c9";
		wait for Clk_period;
		Addr <=  "0010011101110";
		Trees_din <= x"001713c9";
		wait for Clk_period;
		Addr <=  "0010011101111";
		Trees_din <= x"02069e04";
		wait for Clk_period;
		Addr <=  "0010011110000";
		Trees_din <= x"002113c9";
		wait for Clk_period;
		Addr <=  "0010011110001";
		Trees_din <= x"ff5a13c9";
		wait for Clk_period;
		Addr <=  "0010011110010";
		Trees_din <= x"06fedb0c";
		wait for Clk_period;
		Addr <=  "0010011110011";
		Trees_din <= x"01068108";
		wait for Clk_period;
		Addr <=  "0010011110100";
		Trees_din <= x"07026504";
		wait for Clk_period;
		Addr <=  "0010011110101";
		Trees_din <= x"ff971465";
		wait for Clk_period;
		Addr <=  "0010011110110";
		Trees_din <= x"006c1465";
		wait for Clk_period;
		Addr <=  "0010011110111";
		Trees_din <= x"ff721465";
		wait for Clk_period;
		Addr <=  "0010011111000";
		Trees_din <= x"00099624";
		wait for Clk_period;
		Addr <=  "0010011111001";
		Trees_din <= x"010e7620";
		wait for Clk_period;
		Addr <=  "0010011111010";
		Trees_din <= x"0700e910";
		wait for Clk_period;
		Addr <=  "0010011111011";
		Trees_din <= x"02068c08";
		wait for Clk_period;
		Addr <=  "0010011111100";
		Trees_din <= x"05f75104";
		wait for Clk_period;
		Addr <=  "0010011111101";
		Trees_din <= x"00a51465";
		wait for Clk_period;
		Addr <=  "0010011111110";
		Trees_din <= x"00211465";
		wait for Clk_period;
		Addr <=  "0010011111111";
		Trees_din <= x"0c009f04";
		wait for Clk_period;
		Addr <=  "0010100000000";
		Trees_din <= x"ffd41465";
		wait for Clk_period;
		Addr <=  "0010100000001";
		Trees_din <= x"001f1465";
		wait for Clk_period;
		Addr <=  "0010100000010";
		Trees_din <= x"1b026d08";
		wait for Clk_period;
		Addr <=  "0010100000011";
		Trees_din <= x"04fc1d04";
		wait for Clk_period;
		Addr <=  "0010100000100";
		Trees_din <= x"ffef1465";
		wait for Clk_period;
		Addr <=  "0010100000101";
		Trees_din <= x"ff831465";
		wait for Clk_period;
		Addr <=  "0010100000110";
		Trees_din <= x"06058304";
		wait for Clk_period;
		Addr <=  "0010100000111";
		Trees_din <= x"ffc51465";
		wait for Clk_period;
		Addr <=  "0010100001000";
		Trees_din <= x"00571465";
		wait for Clk_period;
		Addr <=  "0010100001001";
		Trees_din <= x"ff871465";
		wait for Clk_period;
		Addr <=  "0010100001010";
		Trees_din <= x"1302970c";
		wait for Clk_period;
		Addr <=  "0010100001011";
		Trees_din <= x"0204ed04";
		wait for Clk_period;
		Addr <=  "0010100001100";
		Trees_din <= x"009e1465";
		wait for Clk_period;
		Addr <=  "0010100001101";
		Trees_din <= x"17faaa04";
		wait for Clk_period;
		Addr <=  "0010100001110";
		Trees_din <= x"ff8e1465";
		wait for Clk_period;
		Addr <=  "0010100001111";
		Trees_din <= x"00781465";
		wait for Clk_period;
		Addr <=  "0010100010000";
		Trees_din <= x"0a003e0c";
		wait for Clk_period;
		Addr <=  "0010100010001";
		Trees_din <= x"0108e508";
		wait for Clk_period;
		Addr <=  "0010100010010";
		Trees_din <= x"08003904";
		wait for Clk_period;
		Addr <=  "0010100010011";
		Trees_din <= x"00651465";
		wait for Clk_period;
		Addr <=  "0010100010100";
		Trees_din <= x"fff01465";
		wait for Clk_period;
		Addr <=  "0010100010101";
		Trees_din <= x"ffa01465";
		wait for Clk_period;
		Addr <=  "0010100010110";
		Trees_din <= x"05f19304";
		wait for Clk_period;
		Addr <=  "0010100010111";
		Trees_din <= x"00031465";
		wait for Clk_period;
		Addr <=  "0010100011000";
		Trees_din <= x"ff6f1465";
		wait for Clk_period;
		Addr <=  "0010100011001";
		Trees_din <= x"010ae22c";
		wait for Clk_period;
		Addr <=  "0010100011010";
		Trees_din <= x"000cd328";
		wait for Clk_period;
		Addr <=  "0010100011011";
		Trees_din <= x"2003ff08";
		wait for Clk_period;
		Addr <=  "0010100011100";
		Trees_din <= x"0b008d04";
		wait for Clk_period;
		Addr <=  "0010100011101";
		Trees_din <= x"ff871509";
		wait for Clk_period;
		Addr <=  "0010100011110";
		Trees_din <= x"ffe11509";
		wait for Clk_period;
		Addr <=  "0010100011111";
		Trees_din <= x"20040010";
		wait for Clk_period;
		Addr <=  "0010100100000";
		Trees_din <= x"08004508";
		wait for Clk_period;
		Addr <=  "0010100100001";
		Trees_din <= x"19000804";
		wait for Clk_period;
		Addr <=  "0010100100010";
		Trees_din <= x"007f1509";
		wait for Clk_period;
		Addr <=  "0010100100011";
		Trees_din <= x"00001509";
		wait for Clk_period;
		Addr <=  "0010100100100";
		Trees_din <= x"1800cd04";
		wait for Clk_period;
		Addr <=  "0010100100101";
		Trees_din <= x"ffa21509";
		wait for Clk_period;
		Addr <=  "0010100100110";
		Trees_din <= x"00191509";
		wait for Clk_period;
		Addr <=  "0010100100111";
		Trees_din <= x"03fa2a08";
		wait for Clk_period;
		Addr <=  "0010100101000";
		Trees_din <= x"08003304";
		wait for Clk_period;
		Addr <=  "0010100101001";
		Trees_din <= x"ffa51509";
		wait for Clk_period;
		Addr <=  "0010100101010";
		Trees_din <= x"001d1509";
		wait for Clk_period;
		Addr <=  "0010100101011";
		Trees_din <= x"0608d704";
		wait for Clk_period;
		Addr <=  "0010100101100";
		Trees_din <= x"ffac1509";
		wait for Clk_period;
		Addr <=  "0010100101101";
		Trees_din <= x"00621509";
		wait for Clk_period;
		Addr <=  "0010100101110";
		Trees_din <= x"ff7f1509";
		wait for Clk_period;
		Addr <=  "0010100101111";
		Trees_din <= x"07fa5b1c";
		wait for Clk_period;
		Addr <=  "0010100110000";
		Trees_din <= x"1b027114";
		wait for Clk_period;
		Addr <=  "0010100110001";
		Trees_din <= x"04ff0d08";
		wait for Clk_period;
		Addr <=  "0010100110010";
		Trees_din <= x"15004704";
		wait for Clk_period;
		Addr <=  "0010100110011";
		Trees_din <= x"001a1509";
		wait for Clk_period;
		Addr <=  "0010100110100";
		Trees_din <= x"00d31509";
		wait for Clk_period;
		Addr <=  "0010100110101";
		Trees_din <= x"0f001404";
		wait for Clk_period;
		Addr <=  "0010100110110";
		Trees_din <= x"ff8a1509";
		wait for Clk_period;
		Addr <=  "0010100110111";
		Trees_din <= x"0a004a04";
		wait for Clk_period;
		Addr <=  "0010100111000";
		Trees_din <= x"00001509";
		wait for Clk_period;
		Addr <=  "0010100111001";
		Trees_din <= x"00951509";
		wait for Clk_period;
		Addr <=  "0010100111010";
		Trees_din <= x"0204b604";
		wait for Clk_period;
		Addr <=  "0010100111011";
		Trees_din <= x"fffe1509";
		wait for Clk_period;
		Addr <=  "0010100111100";
		Trees_din <= x"ff801509";
		wait for Clk_period;
		Addr <=  "0010100111101";
		Trees_din <= x"0f00d704";
		wait for Clk_period;
		Addr <=  "0010100111110";
		Trees_din <= x"ff6f1509";
		wait for Clk_period;
		Addr <=  "0010100111111";
		Trees_din <= x"04fed004";
		wait for Clk_period;
		Addr <=  "0010101000000";
		Trees_din <= x"ffa01509";
		wait for Clk_period;
		Addr <=  "0010101000001";
		Trees_din <= x"00861509";
		wait for Clk_period;
		Addr <=  "0010101000010";
		Trees_din <= x"06ff080c";
		wait for Clk_period;
		Addr <=  "0010101000011";
		Trees_din <= x"1af8f804";
		wait for Clk_period;
		Addr <=  "0010101000100";
		Trees_din <= x"003115a5";
		wait for Clk_period;
		Addr <=  "0010101000101";
		Trees_din <= x"0209d004";
		wait for Clk_period;
		Addr <=  "0010101000110";
		Trees_din <= x"ff7315a5";
		wait for Clk_period;
		Addr <=  "0010101000111";
		Trees_din <= x"002815a5";
		wait for Clk_period;
		Addr <=  "0010101001000";
		Trees_din <= x"00099628";
		wait for Clk_period;
		Addr <=  "0010101001001";
		Trees_din <= x"2003ff08";
		wait for Clk_period;
		Addr <=  "0010101001010";
		Trees_din <= x"0b008d04";
		wait for Clk_period;
		Addr <=  "0010101001011";
		Trees_din <= x"ff8d15a5";
		wait for Clk_period;
		Addr <=  "0010101001100";
		Trees_din <= x"ffe515a5";
		wait for Clk_period;
		Addr <=  "0010101001101";
		Trees_din <= x"20040010";
		wait for Clk_period;
		Addr <=  "0010101001110";
		Trees_din <= x"08004408";
		wait for Clk_period;
		Addr <=  "0010101001111";
		Trees_din <= x"0900e004";
		wait for Clk_period;
		Addr <=  "0010101010000";
		Trees_din <= x"008115a5";
		wait for Clk_period;
		Addr <=  "0010101010001";
		Trees_din <= x"000f15a5";
		wait for Clk_period;
		Addr <=  "0010101010010";
		Trees_din <= x"18020204";
		wait for Clk_period;
		Addr <=  "0010101010011";
		Trees_din <= x"ffa115a5";
		wait for Clk_period;
		Addr <=  "0010101010100";
		Trees_din <= x"003d15a5";
		wait for Clk_period;
		Addr <=  "0010101010101";
		Trees_din <= x"0900d408";
		wait for Clk_period;
		Addr <=  "0010101010110";
		Trees_din <= x"0604ff04";
		wait for Clk_period;
		Addr <=  "0010101010111";
		Trees_din <= x"ff9215a5";
		wait for Clk_period;
		Addr <=  "0010101011000";
		Trees_din <= x"000815a5";
		wait for Clk_period;
		Addr <=  "0010101011001";
		Trees_din <= x"04008e04";
		wait for Clk_period;
		Addr <=  "0010101011010";
		Trees_din <= x"003c15a5";
		wait for Clk_period;
		Addr <=  "0010101011011";
		Trees_din <= x"ffcb15a5";
		wait for Clk_period;
		Addr <=  "0010101011100";
		Trees_din <= x"08004c18";
		wait for Clk_period;
		Addr <=  "0010101011101";
		Trees_din <= x"0401ac08";
		wait for Clk_period;
		Addr <=  "0010101011110";
		Trees_din <= x"1c028404";
		wait for Clk_period;
		Addr <=  "0010101011111";
		Trees_din <= x"ff7215a5";
		wait for Clk_period;
		Addr <=  "0010101100000";
		Trees_din <= x"ffe715a5";
		wait for Clk_period;
		Addr <=  "0010101100001";
		Trees_din <= x"000b8f08";
		wait for Clk_period;
		Addr <=  "0010101100010";
		Trees_din <= x"02044d04";
		wait for Clk_period;
		Addr <=  "0010101100011";
		Trees_din <= x"008a15a5";
		wait for Clk_period;
		Addr <=  "0010101100100";
		Trees_din <= x"001915a5";
		wait for Clk_period;
		Addr <=  "0010101100101";
		Trees_din <= x"03f4de04";
		wait for Clk_period;
		Addr <=  "0010101100110";
		Trees_din <= x"000515a5";
		wait for Clk_period;
		Addr <=  "0010101100111";
		Trees_din <= x"ff9215a5";
		wait for Clk_period;
		Addr <=  "0010101101000";
		Trees_din <= x"007f15a5";
		wait for Clk_period;
		Addr <=  "0010101101001";
		Trees_din <= x"0604df40";
		wait for Clk_period;
		Addr <=  "0010101101010";
		Trees_din <= x"00036a08";
		wait for Clk_period;
		Addr <=  "0010101101011";
		Trees_din <= x"0c007604";
		wait for Clk_period;
		Addr <=  "0010101101100";
		Trees_din <= x"002a16b9";
		wait for Clk_period;
		Addr <=  "0010101101101";
		Trees_din <= x"ff6e16b9";
		wait for Clk_period;
		Addr <=  "0010101101110";
		Trees_din <= x"0006361c";
		wait for Clk_period;
		Addr <=  "0010101101111";
		Trees_din <= x"0104940c";
		wait for Clk_period;
		Addr <=  "0010101110000";
		Trees_din <= x"11013904";
		wait for Clk_period;
		Addr <=  "0010101110001";
		Trees_din <= x"00ea16b9";
		wait for Clk_period;
		Addr <=  "0010101110010";
		Trees_din <= x"0d00a304";
		wait for Clk_period;
		Addr <=  "0010101110011";
		Trees_din <= x"005416b9";
		wait for Clk_period;
		Addr <=  "0010101110100";
		Trees_din <= x"ffa716b9";
		wait for Clk_period;
		Addr <=  "0010101110101";
		Trees_din <= x"0b007008";
		wait for Clk_period;
		Addr <=  "0010101110110";
		Trees_din <= x"0b006d04";
		wait for Clk_period;
		Addr <=  "0010101110111";
		Trees_din <= x"ffcb16b9";
		wait for Clk_period;
		Addr <=  "0010101111000";
		Trees_din <= x"00d116b9";
		wait for Clk_period;
		Addr <=  "0010101111001";
		Trees_din <= x"11027504";
		wait for Clk_period;
		Addr <=  "0010101111010";
		Trees_din <= x"ff8016b9";
		wait for Clk_period;
		Addr <=  "0010101111011";
		Trees_din <= x"004116b9";
		wait for Clk_period;
		Addr <=  "0010101111100";
		Trees_din <= x"03fab210";
		wait for Clk_period;
		Addr <=  "0010101111101";
		Trees_din <= x"09009408";
		wait for Clk_period;
		Addr <=  "0010101111110";
		Trees_din <= x"1f027604";
		wait for Clk_period;
		Addr <=  "0010101111111";
		Trees_din <= x"007116b9";
		wait for Clk_period;
		Addr <=  "0010110000000";
		Trees_din <= x"ff9216b9";
		wait for Clk_period;
		Addr <=  "0010110000001";
		Trees_din <= x"0f015704";
		wait for Clk_period;
		Addr <=  "0010110000010";
		Trees_din <= x"ff7f16b9";
		wait for Clk_period;
		Addr <=  "0010110000011";
		Trees_din <= x"001f16b9";
		wait for Clk_period;
		Addr <=  "0010110000100";
		Trees_din <= x"0b006908";
		wait for Clk_period;
		Addr <=  "0010110000101";
		Trees_din <= x"0b006404";
		wait for Clk_period;
		Addr <=  "0010110000110";
		Trees_din <= x"001716b9";
		wait for Clk_period;
		Addr <=  "0010110000111";
		Trees_din <= x"00ae16b9";
		wait for Clk_period;
		Addr <=  "0010110001000";
		Trees_din <= x"ffb216b9";
		wait for Clk_period;
		Addr <=  "0010110001001";
		Trees_din <= x"0106182c";
		wait for Clk_period;
		Addr <=  "0010110001010";
		Trees_din <= x"0607fa14";
		wait for Clk_period;
		Addr <=  "0010110001011";
		Trees_din <= x"0207e90c";
		wait for Clk_period;
		Addr <=  "0010110001100";
		Trees_din <= x"17f75604";
		wait for Clk_period;
		Addr <=  "0010110001101";
		Trees_din <= x"006516b9";
		wait for Clk_period;
		Addr <=  "0010110001110";
		Trees_din <= x"1afc4504";
		wait for Clk_period;
		Addr <=  "0010110001111";
		Trees_din <= x"002416b9";
		wait for Clk_period;
		Addr <=  "0010110010000";
		Trees_din <= x"ff8016b9";
		wait for Clk_period;
		Addr <=  "0010110010001";
		Trees_din <= x"1b025104";
		wait for Clk_period;
		Addr <=  "0010110010010";
		Trees_din <= x"fffd16b9";
		wait for Clk_period;
		Addr <=  "0010110010011";
		Trees_din <= x"ff7216b9";
		wait for Clk_period;
		Addr <=  "0010110010100";
		Trees_din <= x"15004810";
		wait for Clk_period;
		Addr <=  "0010110010101";
		Trees_din <= x"15003f08";
		wait for Clk_period;
		Addr <=  "0010110010110";
		Trees_din <= x"03f80c04";
		wait for Clk_period;
		Addr <=  "0010110010111";
		Trees_din <= x"000116b9";
		wait for Clk_period;
		Addr <=  "0010110011000";
		Trees_din <= x"007516b9";
		wait for Clk_period;
		Addr <=  "0010110011001";
		Trees_din <= x"11024404";
		wait for Clk_period;
		Addr <=  "0010110011010";
		Trees_din <= x"ff9316b9";
		wait for Clk_period;
		Addr <=  "0010110011011";
		Trees_din <= x"006416b9";
		wait for Clk_period;
		Addr <=  "0010110011100";
		Trees_din <= x"04013604";
		wait for Clk_period;
		Addr <=  "0010110011101";
		Trees_din <= x"008716b9";
		wait for Clk_period;
		Addr <=  "0010110011110";
		Trees_din <= x"fff916b9";
		wait for Clk_period;
		Addr <=  "0010110011111";
		Trees_din <= x"0f00030c";
		wait for Clk_period;
		Addr <=  "0010110100000";
		Trees_din <= x"02066208";
		wait for Clk_period;
		Addr <=  "0010110100001";
		Trees_din <= x"04fc2904";
		wait for Clk_period;
		Addr <=  "0010110100010";
		Trees_din <= x"ffdc16b9";
		wait for Clk_period;
		Addr <=  "0010110100011";
		Trees_din <= x"004516b9";
		wait for Clk_period;
		Addr <=  "0010110100100";
		Trees_din <= x"ff8616b9";
		wait for Clk_period;
		Addr <=  "0010110100101";
		Trees_din <= x"03fa1410";
		wait for Clk_period;
		Addr <=  "0010110100110";
		Trees_din <= x"03f5db08";
		wait for Clk_period;
		Addr <=  "0010110100111";
		Trees_din <= x"0a004104";
		wait for Clk_period;
		Addr <=  "0010110101000";
		Trees_din <= x"002816b9";
		wait for Clk_period;
		Addr <=  "0010110101001";
		Trees_din <= x"ffcc16b9";
		wait for Clk_period;
		Addr <=  "0010110101010";
		Trees_din <= x"04fc2904";
		wait for Clk_period;
		Addr <=  "0010110101011";
		Trees_din <= x"000116b9";
		wait for Clk_period;
		Addr <=  "0010110101100";
		Trees_din <= x"00a616b9";
		wait for Clk_period;
		Addr <=  "0010110101101";
		Trees_din <= x"ffca16b9";
		wait for Clk_period;
		Addr <=  "0010110101110";
		Trees_din <= x"010ae23c";
		wait for Clk_period;
		Addr <=  "0010110101111";
		Trees_din <= x"000cd338";
		wait for Clk_period;
		Addr <=  "0010110110000";
		Trees_din <= x"00034418";
		wait for Clk_period;
		Addr <=  "0010110110001";
		Trees_din <= x"06058308";
		wait for Clk_period;
		Addr <=  "0010110110010";
		Trees_din <= x"12006204";
		wait for Clk_period;
		Addr <=  "0010110110011";
		Trees_din <= x"0027176d";
		wait for Clk_period;
		Addr <=  "0010110110100";
		Trees_din <= x"ff78176d";
		wait for Clk_period;
		Addr <=  "0010110110101";
		Trees_din <= x"11001008";
		wait for Clk_period;
		Addr <=  "0010110110110";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0010110110111";
		Trees_din <= x"ffe4176d";
		wait for Clk_period;
		Addr <=  "0010110111000";
		Trees_din <= x"ff88176d";
		wait for Clk_period;
		Addr <=  "0010110111001";
		Trees_din <= x"15004804";
		wait for Clk_period;
		Addr <=  "0010110111010";
		Trees_din <= x"000d176d";
		wait for Clk_period;
		Addr <=  "0010110111011";
		Trees_din <= x"0077176d";
		wait for Clk_period;
		Addr <=  "0010110111100";
		Trees_din <= x"0c009c10";
		wait for Clk_period;
		Addr <=  "0010110111101";
		Trees_din <= x"1b024508";
		wait for Clk_period;
		Addr <=  "0010110111110";
		Trees_din <= x"0d000f04";
		wait for Clk_period;
		Addr <=  "0010110111111";
		Trees_din <= x"000a176d";
		wait for Clk_period;
		Addr <=  "0010111000000";
		Trees_din <= x"008f176d";
		wait for Clk_period;
		Addr <=  "0010111000001";
		Trees_din <= x"0e004504";
		wait for Clk_period;
		Addr <=  "0010111000010";
		Trees_din <= x"ff9c176d";
		wait for Clk_period;
		Addr <=  "0010111000011";
		Trees_din <= x"0024176d";
		wait for Clk_period;
		Addr <=  "0010111000100";
		Trees_din <= x"00077208";
		wait for Clk_period;
		Addr <=  "0010111000101";
		Trees_din <= x"0a003e04";
		wait for Clk_period;
		Addr <=  "0010111000110";
		Trees_din <= x"ffe5176d";
		wait for Clk_period;
		Addr <=  "0010111000111";
		Trees_din <= x"0064176d";
		wait for Clk_period;
		Addr <=  "0010111001000";
		Trees_din <= x"11020604";
		wait for Clk_period;
		Addr <=  "0010111001001";
		Trees_din <= x"ffc9176d";
		wait for Clk_period;
		Addr <=  "0010111001010";
		Trees_din <= x"004b176d";
		wait for Clk_period;
		Addr <=  "0010111001011";
		Trees_din <= x"ff89176d";
		wait for Clk_period;
		Addr <=  "0010111001100";
		Trees_din <= x"04fe9608";
		wait for Clk_period;
		Addr <=  "0010111001101";
		Trees_din <= x"10005604";
		wait for Clk_period;
		Addr <=  "0010111001110";
		Trees_din <= x"ff73176d";
		wait for Clk_period;
		Addr <=  "0010111001111";
		Trees_din <= x"0030176d";
		wait for Clk_period;
		Addr <=  "0010111010000";
		Trees_din <= x"04ff0d08";
		wait for Clk_period;
		Addr <=  "0010111010001";
		Trees_din <= x"1101f004";
		wait for Clk_period;
		Addr <=  "0010111010010";
		Trees_din <= x"0011176d";
		wait for Clk_period;
		Addr <=  "0010111010011";
		Trees_din <= x"00c8176d";
		wait for Clk_period;
		Addr <=  "0010111010100";
		Trees_din <= x"0604df08";
		wait for Clk_period;
		Addr <=  "0010111010101";
		Trees_din <= x"1402bc04";
		wait for Clk_period;
		Addr <=  "0010111010110";
		Trees_din <= x"002c176d";
		wait for Clk_period;
		Addr <=  "0010111010111";
		Trees_din <= x"ff7a176d";
		wait for Clk_period;
		Addr <=  "0010111011000";
		Trees_din <= x"03f7de04";
		wait for Clk_period;
		Addr <=  "0010111011001";
		Trees_din <= x"fff5176d";
		wait for Clk_period;
		Addr <=  "0010111011010";
		Trees_din <= x"0072176d";
		wait for Clk_period;
		Addr <=  "0010111011011";
		Trees_din <= x"06fedb0c";
		wait for Clk_period;
		Addr <=  "0010111011100";
		Trees_din <= x"01068108";
		wait for Clk_period;
		Addr <=  "0010111011101";
		Trees_din <= x"05f6ed04";
		wait for Clk_period;
		Addr <=  "0010111011110";
		Trees_din <= x"00671819";
		wait for Clk_period;
		Addr <=  "0010111011111";
		Trees_din <= x"ffaa1819";
		wait for Clk_period;
		Addr <=  "0010111100000";
		Trees_din <= x"ff7b1819";
		wait for Clk_period;
		Addr <=  "0010111100001";
		Trees_din <= x"0700e934";
		wait for Clk_period;
		Addr <=  "0010111100010";
		Trees_din <= x"02050518";
		wait for Clk_period;
		Addr <=  "0010111100011";
		Trees_din <= x"0a004810";
		wait for Clk_period;
		Addr <=  "0010111100100";
		Trees_din <= x"19000908";
		wait for Clk_period;
		Addr <=  "0010111100101";
		Trees_din <= x"0b005a04";
		wait for Clk_period;
		Addr <=  "0010111100110";
		Trees_din <= x"ffc11819";
		wait for Clk_period;
		Addr <=  "0010111100111";
		Trees_din <= x"00851819";
		wait for Clk_period;
		Addr <=  "0010111101000";
		Trees_din <= x"07fc8f04";
		wait for Clk_period;
		Addr <=  "0010111101001";
		Trees_din <= x"00181819";
		wait for Clk_period;
		Addr <=  "0010111101010";
		Trees_din <= x"ffa91819";
		wait for Clk_period;
		Addr <=  "0010111101011";
		Trees_din <= x"0604df04";
		wait for Clk_period;
		Addr <=  "0010111101100";
		Trees_din <= x"ff991819";
		wait for Clk_period;
		Addr <=  "0010111101101";
		Trees_din <= x"002e1819";
		wait for Clk_period;
		Addr <=  "0010111101110";
		Trees_din <= x"0605ab0c";
		wait for Clk_period;
		Addr <=  "0010111101111";
		Trees_din <= x"05f40e04";
		wait for Clk_period;
		Addr <=  "0010111110000";
		Trees_din <= x"ff821819";
		wait for Clk_period;
		Addr <=  "0010111110001";
		Trees_din <= x"0b009f04";
		wait for Clk_period;
		Addr <=  "0010111110010";
		Trees_din <= x"ffe31819";
		wait for Clk_period;
		Addr <=  "0010111110011";
		Trees_din <= x"00681819";
		wait for Clk_period;
		Addr <=  "0010111110100";
		Trees_din <= x"07fbe808";
		wait for Clk_period;
		Addr <=  "0010111110101";
		Trees_din <= x"0007d404";
		wait for Clk_period;
		Addr <=  "0010111110110";
		Trees_din <= x"004f1819";
		wait for Clk_period;
		Addr <=  "0010111110111";
		Trees_din <= x"ffbb1819";
		wait for Clk_period;
		Addr <=  "0010111111000";
		Trees_din <= x"0e002e04";
		wait for Clk_period;
		Addr <=  "0010111111001";
		Trees_din <= x"00291819";
		wait for Clk_period;
		Addr <=  "0010111111010";
		Trees_din <= x"ffbe1819";
		wait for Clk_period;
		Addr <=  "0010111111011";
		Trees_din <= x"1b026d08";
		wait for Clk_period;
		Addr <=  "0010111111100";
		Trees_din <= x"04fc1d04";
		wait for Clk_period;
		Addr <=  "0010111111101";
		Trees_din <= x"ffe41819";
		wait for Clk_period;
		Addr <=  "0010111111110";
		Trees_din <= x"ff871819";
		wait for Clk_period;
		Addr <=  "0010111111111";
		Trees_din <= x"06058308";
		wait for Clk_period;
		Addr <=  "0011000000000";
		Trees_din <= x"01000504";
		wait for Clk_period;
		Addr <=  "0011000000001";
		Trees_din <= x"00301819";
		wait for Clk_period;
		Addr <=  "0011000000010";
		Trees_din <= x"ff981819";
		wait for Clk_period;
		Addr <=  "0011000000011";
		Trees_din <= x"05f95b04";
		wait for Clk_period;
		Addr <=  "0011000000100";
		Trees_din <= x"00721819";
		wait for Clk_period;
		Addr <=  "0011000000101";
		Trees_din <= x"ffe31819";
		wait for Clk_period;
		Addr <=  "0011000000110";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  5
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"04080d64";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"04039038";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"1c02871c";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"0400170c";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"0c003f08";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"010a5104";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"ff900105";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"00370105";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"ff540105";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"0d000008";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"0c009704";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"ff700105";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"00590105";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"05f55604";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"ff560105";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"ff7a0105";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"04ffbc0c";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"0b006608";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"00061604";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"00370105";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"ffa40105";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"ff580105";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"12007808";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"03f4de04";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"00370105";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"ff790105";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"0c00c204";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"019a0105";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"ff8c0105";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"000d411c";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"020ab010";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"03f6c208";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"15003404";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"00ca0105";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"ff740105";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"06fe5904";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"001e0105";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"02760105";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"16006308";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"0b007504";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"012b0105";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"ff7e0105";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"ff600105";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"1103010c";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"08004b04";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"ff540105";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"01054b04";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"ff8c0105";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"00370105";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"000f0105";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"00120e18";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"020d7910";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"0109880c";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"15004c08";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"08003604";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"012b0105";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"03c20105";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"00370105";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"ff900105";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"11009604";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"00ca0105";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"ff840105";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"07fc0d04";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"ff5e0105";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"00370105";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"0403e740";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"1c028728";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"0400170c";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"0c003f08";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"11000004";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"00430201";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"ff9a0201";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"ff5a0201";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"07ff330c";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"1cfd6d04";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"00170201";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"0d000004";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"ffa70201";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"ff680201";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"11002608";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"0f000104";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"00050201";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"016c0201";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"04039004";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"ff750201";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"00e50201";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"04ffbc08";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"17f98104";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"fff60201";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"ff5f0201";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"0e00350c";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"0c00b104";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"ff760201";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"10003e04";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"ff840201";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"01680201";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"01440201";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"000d411c";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"020d7914";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"010dc810";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"04057d08";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"020ab004";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"013f0201";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"ff7e0201";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"0109ed04";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"02070201";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"ff9e0201";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"ff8a0201";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"08004504";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"ff6a0201";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"00320201";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"040a8414";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"13021808";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"1301b404";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"ff7e0201";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"00fe0201";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"08004b04";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"ff5a0201";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"0a004f04";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"ffa30201";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"003a0201";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"0010df08";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"05f80604";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"017e0201";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"000e0201";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"0f019904";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"ff760201";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"00410201";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"0403e740";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"1c028728";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"0400170c";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"0b004708";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"0a003804";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"004302d5";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"ff9f02d5";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"ff5f02d5";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"07ff330c";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"1cfd6d04";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"001602d5";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"04002b04";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"ffde02d5";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"ff7102d5";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"0208b708";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"0f001e04";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"ff6902d5";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"002502d5";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"07ff8f04";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"016b02d5";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"000302d5";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"04ffbc08";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"0b006604";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"000302d5";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"ff6402d5";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"02076e0c";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"16005b04";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"ff8d02d5";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"1d028804";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"015802d5";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"ff9a02d5";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"ff8702d5";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"0010df24";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"020d791c";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"0109ed10";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"04057d08";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"1b028304";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"000302d5";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"015202d5";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"18000a04";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"004a02d5";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"014f02d5";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"17f72e04";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"011002d5";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"08004504";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"ff6902d5";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"008302d5";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"08004804";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"ff6a02d5";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"008e02d5";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"10003004";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"008602d5";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"ff5e02d5";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"0403e73c";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"04ffbc08";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"17f69904";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"fff903c9";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"ff6303c9";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"1c028720";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"07ff3310";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"05f54508";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"0d000004";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"ffbc03c9";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"ff6503c9";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"05f55d04";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"005f03c9";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"ff8b03c9";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"0208e008";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"04039004";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"ff8e03c9";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"008303c9";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"11002604";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"015e03c9";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"ffe803c9";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"0e00350c";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"0c00b104";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"ff7d03c9";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"10003e04";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"ff9103c9";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"00df03c9";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"02045404";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"015303c9";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"002603c9";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"000d4120";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"020d7918";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"16005308";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"10003404";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"002003c9";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"ff8003c9";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"0b006508";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"17f75c04";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"00d503c9";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"ff7503c9";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"0d000a04";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"005b03c9";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"012f03c9";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"08004804";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"ff7503c9";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"003803c9";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"040a8410";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"13021808";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"1301b404";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"ff8b03c9";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"00d003c9";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"08004b04";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"ff6103c9";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"fff903c9";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"07fb4d0c";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"0a005008";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"0107ce04";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"ff7103c9";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"002003c9";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"00d003c9";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"014103c9";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"04032340";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"1c028724";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"04001708";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"0c003f04";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"000604a5";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"ff6604a5";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"07fb190c";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"1e061a08";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"04001f04";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"002304a5";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"ff6804a5";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"002a04a5";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"0c00a108";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"0e004c04";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"ff6604a5";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"ffef04a5";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"0c00a704";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"013d04a5";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"ffa904a5";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"04ffbc08";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"17f98104";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"002704a5";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"ff6c04a5";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"0e003510";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"0e002808";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"1f028804";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"fffc04a5";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"00d704a5";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"09007804";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"002d04a5";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"ff7c04a5";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"00f904a5";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"000e8018";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"020f5a14";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"010dc810";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"16005308";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"0602d004";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"ff7b04a5";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"002104a5";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"02076e04";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"00fa04a5";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"006a04a5";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"ff7d04a5";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"ff7804a5";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"0408b408";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"22000004";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"ff6304a5";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"003b04a5";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"03f51804";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"ff7d04a5";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"18001b04";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"ff9304a5";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"05f59704";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"fffa04a5";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"00f804a5";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"04032340";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"1c028728";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"04001708";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"0e005c04";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"ff690591";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"000d0591";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"07fb1910";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"0d000008";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"08004204";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"ff820591";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"00c20591";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"1e061a04";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"ff670591";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"003f0591";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"0c00a108";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"0e004c04";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"ff6a0591";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"fff40591";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"0c00a704";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"00e90591";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"ffb30591";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"04ffbc08";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"0b006604";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"00300591";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"ff710591";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"0110a10c";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"010d0c08";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"05f7db04";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"ff850591";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"00920591";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"010b0591";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"ff9b0591";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"0010df30";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"07fb5f1c";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"0408b410";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"06feca08";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"0e003104";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"ffca0591";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"01230591";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"09007004";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"008c0591";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"ffa80591";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"08002d04";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"ff9c0591";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"0f00bc04";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"00cc0591";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"ffec0591";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"01f5d104";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"ff920591";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"03f7b908";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"0d002304";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"ff940591";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"007a0591";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"09009704";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"00710591";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"01260591";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"0c010904";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"ff670591";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"00770591";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"04032340";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"1c028724";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"04ffdd08";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"17f69904";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"00190665";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"ff6c0665";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"0d00000c";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"0c009704";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"ff790665";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"1afb7a04";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"01a80665";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"00030665";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"05f54508";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"04002b04";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"ffa30665";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"ff650665";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"01084c04";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"ff860665";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"fff20665";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"04ffbc08";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"17f98104";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"003a0665";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"ff750665";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"1d028810";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"0a003f08";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"08003e04";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"ff9b0665";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"00310665";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"0f009404";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"00030665";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"00f00665";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"ff9f0665";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"0010df24";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"010dc820";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"020ab010";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"10004808";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"0d007f04";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"ffab0665";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"009d0665";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"05f4f804";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"001f0665";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"00dc0665";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"04098208";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"16006304";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"000e0665";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"ff690665";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"0f000404";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"ffdb0665";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"00c80665";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"ff7c0665";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"0c010904";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"ff6a0665";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"006c0665";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"0403233c";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"1c028724";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"04ffdd08";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"0c003f04";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"00230771";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"ff6f0771";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"010b6e10";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"0d000208";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"1afcea04";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"00c10771";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"ff920771";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"01084c04";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"ff870771";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"fffb0771";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"0f000308";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"0c00b004";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"ff720771";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"00850771";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"ff670771";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"04ffbc08";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"0b006604";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"003d0771";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"ff790771";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"0900e50c";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"16005b04";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"ffa40771";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"02069e04";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"00d80771";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"ffef0771";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"ffa30771";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"000e8034";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"0a004114";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"0e002f08";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"1f025804";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"001f0771";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"ff660771";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"0205ff04";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"00e30771";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"03f91804";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"ff940771";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"00710771";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"03f7ad10";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"04067d08";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"15003404";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"00710771";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"ff900771";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"0d000804";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"ff970771";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"00ae0771";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"03fa0a08";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"0e002304";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"ffe60771";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"00d40771";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"0a004604";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"00890771";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"ffc30771";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"0408b408";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"19004f04";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"ff6a0771";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"00310771";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"0800420c";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"020ab008";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"07f8a004";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"fff70771";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"00c80771";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"ffa60771";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"ff860771";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"04032344";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"04ff7c14";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"17f69904";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"00370865";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"0d008d04";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"ff640865";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"0d009504";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"006d0865";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"11009a04";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"002d0865";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"ff7a0865";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"0900b818";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"0900a60c";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"02030504";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"00ad0865";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"06fd7604";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"003c0865";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"ff8c0865";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"07f91e04";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"ff8d0865";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"1c025704";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"ff9d0865";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"01520865";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"1c028810";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"1102dd08";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"03fb2d04";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"ff700865";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"00280865";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"05f55604";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"ffa90865";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"00db0865";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"0c00b104";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"ff970865";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"00ad0865";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"0010df30";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"07fb5f1c";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"1302570c";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"020b0308";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"000c8b04";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"00530865";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"01280865";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"ffa50865";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"1b026608";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"18000004";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"009f0865";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"ff870865";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"0f00bc04";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"00490865";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"ff970865";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"01f5d104";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"ffa50865";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"03f7b908";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"17f82b04";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"00630865";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"ff910865";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"0b006604";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"002c0865";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"00cf0865";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"12009904";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"ff700865";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"005b0865";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"0401f43c";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"04ff7c14";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"0e005c10";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"0d008d04";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"ff650965";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"0d009504";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"00640965";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"11009a04";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"002e0965";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"ff7f0965";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"003e0965";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"0d000510";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"1f025904";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"ff830965";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"08003204";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"ffa80965";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"1b027c04";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"010b0965";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"fffb0965";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"0206b910";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"0205c008";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"1afb5304";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"fff80965";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"ff6c0965";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"0f000c04";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"00d20965";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"ffbb0965";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"03fb4204";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"ff680965";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"00200965";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"05f4fd1c";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"03f89b10";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"06048d08";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"06fcd304";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"fff40965";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"ff670965";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"07f66c04";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"008d0965";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"ff9f0965";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"0b007c08";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"0a004004";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"fff70965";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"ffa40965";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"00a30965";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"03f51808";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"00098404";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"001a0965";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"ff770965";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"08004110";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"04051908";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"1c028004";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"ff930965";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"004c0965";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"05f7a704";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"ffe70965";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"009a0965";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"16007a08";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"0b006604";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"fff40965";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"00da0965";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"0d000104";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"00b20965";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"ffd20965";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"04006334";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"06ff0810";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"1d02880c";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"1102d804";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"ff660a71";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"1c027304";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"004a0a71";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"ff8b0a71";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"fff70a71";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"11000008";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"0006db04";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"ffab0a71";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"00bd0a71";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"07029710";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"06ff2a08";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"0e003104";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"ffa60a71";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"00960a71";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"18000204";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"00090a71";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"ff7a0a71";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"02038904";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"ff820a71";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"0d008a04";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"ffa20a71";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"01290a71";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"05f4fd20";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"0900eb14";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"0408b40c";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"00068c04";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"00340a71";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"1f028804";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"ff670a71";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"002d0a71";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"0e004204";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"ffdc0a71";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"007a0a71";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"10004508";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"0c00a004";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"016b0a71";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"ffac0a71";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"ff880a71";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"13025718";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"13018a08";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"07f93504";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"fff70a71";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"ff990a71";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"06ff6f08";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"0e003a04";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"01500a71";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"00220a71";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"04041d04";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"ffd90a71";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"00890a71";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"07fb3610";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"1e024a08";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"06003004";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"00be0a71";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"ffa00a71";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"04063004";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"ff920a71";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"002f0a71";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"1302ff04";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"ff900a71";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"07ff4304";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"00730a71";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"ffe40a71";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"04ffbc20";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"0b006610";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"16006a04";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"01260b5d";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"08003c08";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"06003f04";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"ff9a0b5d";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"00d10b5d";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"ff6f0b5d";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"0f00020c";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"10004208";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"1100b004";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"ffae0b5d";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"01750b5d";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"ff740b5d";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"ff6b0b5d";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"0900b828";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"000fee1c";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"03f9c510";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"0c00da08";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"0f000104";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"ffe70b5d";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"00950b5d";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"1100d204";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"ffe80b5d";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"ff9b0b5d";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"0403e704";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"ff7d0b5d";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"06ff2a04";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"003a0b5d";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"fff20b5d";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"10003004";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"005e0b5d";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"0f013604";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"ff760b5d";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"00080b5d";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"05f7ca18";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"03fb4210";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"18000008";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"0d000004";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"ffa40b5d";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"00b00b5d";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"13025704";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"00070b5d";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"ff8a0b5d";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"0d003a04";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"000f0b5d";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"00d60b5d";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"0401c208";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"1afa6704";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"00090b5d";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"ff7d0b5d";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"000b6a08";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"01fc5404";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"ffa70b5d";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"00930b5d";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"17f70f04";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"00590b5d";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"ffb50b5d";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"04ffbc28";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"0b006610";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"16006a04";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"00e80c61";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"08003c08";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"06003f04";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"ff9f0c61";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"00b20c61";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"ff710c61";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"0f00020c";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"10004208";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"0a004804";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"ffac0c61";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"013c0c61";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"ff760c61";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"16004e08";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"0b008204";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"00470c61";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"ff7e0c61";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"ff670c61";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"0900b828";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"000ed01c";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"000d8e10";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"04043008";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"07fb1904";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"ff870c61";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"00330c61";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"17f7a404";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"000b0c61";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"00a10c61";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"0a004604";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"fff90c61";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"04020704";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"01b90c61";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"00860c61";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"19002c08";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"040a8404";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"ff770c61";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"00230c61";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"00660c61";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"0402ab18";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"13022b08";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"0900de04";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"ffa00c61";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"00c30c61";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"00123208";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"03fb4204";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"ff710c61";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"00210c61";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"19000104";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"ffae0c61";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"00c20c61";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"000cd30c";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"000c8b08";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"05f77a04";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"ffc10c61";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"005f0c61";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"01220c61";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"0408b408";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"07fc7104";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"ff730c61";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"ffdf0c61";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"06009a04";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"00660c61";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"ffa20c61";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"04ffbc28";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"0b006610";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"0e003508";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"13037e04";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"013a0d6d";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"ff9a0d6d";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"11000004";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"00330d6d";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"ff730d6d";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"0f00020c";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"10004208";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"1100b004";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"ffb00d6d";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"00fe0d6d";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"ff7a0d6d";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"16004e08";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"03fc4004";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"ff810d6d";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"00440d6d";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"ff680d6d";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"0900b834";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"0900ad20";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"0b007c10";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"04080d08";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"19000b04";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"ff720d6d";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"00290d6d";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"000cb204";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"00780d6d";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"00030d6d";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"00088d08";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"11004c04";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"003f0d6d";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"ff850d6d";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"05f57804";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"ffe00d6d";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"00ad0d6d";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"0e003208";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"07fa3c04";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"ff9b0d6d";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"00120d6d";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"0205a804";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"00150d6d";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"0206e604";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"01550d6d";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"006f0d6d";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"03fb2d20";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"05f7ca10";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"0c00a008";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"10004504";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"00aa0d6d";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"ffc10d6d";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"13025704";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"00400d6d";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"ff730d6d";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"0d008208";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"08003804";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"00420d6d";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"ff9a0d6d";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"03f91804";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"00080d6d";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"008c0d6d";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"15003d08";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"0600c004";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"003a0d6d";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"01020d6d";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"ffbc0d6d";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"04ff7c28";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"0b006614";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"16006a08";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"17f7d904";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"00dc0e79";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"00270e79";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"08003c08";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"04fe0304";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"ffa60e79";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"00b50e79";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"ff760e79";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"0f000008";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"11011e04";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"ff890e79";
		wait for Clk_period;
		Addr <=  "0001101101001";
		Trees_din <= x"00d80e79";
		wait for Clk_period;
		Addr <=  "0001101101010";
		Trees_din <= x"16004e08";
		wait for Clk_period;
		Addr <=  "0001101101011";
		Trees_din <= x"0b008204";
		wait for Clk_period;
		Addr <=  "0001101101100";
		Trees_din <= x"00460e79";
		wait for Clk_period;
		Addr <=  "0001101101101";
		Trees_din <= x"ff850e79";
		wait for Clk_period;
		Addr <=  "0001101101110";
		Trees_din <= x"ff690e79";
		wait for Clk_period;
		Addr <=  "0001101101111";
		Trees_din <= x"0900b830";
		wait for Clk_period;
		Addr <=  "0001101110000";
		Trees_din <= x"0900ad1c";
		wait for Clk_period;
		Addr <=  "0001101110001";
		Trees_din <= x"04045610";
		wait for Clk_period;
		Addr <=  "0001101110010";
		Trees_din <= x"06ff2a08";
		wait for Clk_period;
		Addr <=  "0001101110011";
		Trees_din <= x"05f57d04";
		wait for Clk_period;
		Addr <=  "0001101110100";
		Trees_din <= x"ffaa0e79";
		wait for Clk_period;
		Addr <=  "0001101110101";
		Trees_din <= x"009c0e79";
		wait for Clk_period;
		Addr <=  "0001101110110";
		Trees_din <= x"0d000004";
		wait for Clk_period;
		Addr <=  "0001101110111";
		Trees_din <= x"004b0e79";
		wait for Clk_period;
		Addr <=  "0001101111000";
		Trees_din <= x"ff7a0e79";
		wait for Clk_period;
		Addr <=  "0001101111001";
		Trees_din <= x"000fee08";
		wait for Clk_period;
		Addr <=  "0001101111010";
		Trees_din <= x"020b0304";
		wait for Clk_period;
		Addr <=  "0001101111011";
		Trees_din <= x"008e0e79";
		wait for Clk_period;
		Addr <=  "0001101111100";
		Trees_din <= x"fff20e79";
		wait for Clk_period;
		Addr <=  "0001101111101";
		Trees_din <= x"ffbd0e79";
		wait for Clk_period;
		Addr <=  "0001101111110";
		Trees_din <= x"07f91e08";
		wait for Clk_period;
		Addr <=  "0001101111111";
		Trees_din <= x"03f89b04";
		wait for Clk_period;
		Addr <=  "0001110000000";
		Trees_din <= x"ffa30e79";
		wait for Clk_period;
		Addr <=  "0001110000001";
		Trees_din <= x"00350e79";
		wait for Clk_period;
		Addr <=  "0001110000010";
		Trees_din <= x"04002b04";
		wait for Clk_period;
		Addr <=  "0001110000011";
		Trees_din <= x"01420e79";
		wait for Clk_period;
		Addr <=  "0001110000100";
		Trees_din <= x"00086304";
		wait for Clk_period;
		Addr <=  "0001110000101";
		Trees_din <= x"00980e79";
		wait for Clk_period;
		Addr <=  "0001110000110";
		Trees_din <= x"00090e79";
		wait for Clk_period;
		Addr <=  "0001110000111";
		Trees_din <= x"0402ab14";
		wait for Clk_period;
		Addr <=  "0001110001000";
		Trees_din <= x"0900e004";
		wait for Clk_period;
		Addr <=  "0001110001001";
		Trees_din <= x"ff700e79";
		wait for Clk_period;
		Addr <=  "0001110001010";
		Trees_din <= x"10004208";
		wait for Clk_period;
		Addr <=  "0001110001011";
		Trees_din <= x"15003704";
		wait for Clk_period;
		Addr <=  "0001110001100";
		Trees_din <= x"ff9a0e79";
		wait for Clk_period;
		Addr <=  "0001110001101";
		Trees_din <= x"00a50e79";
		wait for Clk_period;
		Addr <=  "0001110001110";
		Trees_din <= x"1c024e04";
		wait for Clk_period;
		Addr <=  "0001110001111";
		Trees_din <= x"00180e79";
		wait for Clk_period;
		Addr <=  "0001110010000";
		Trees_din <= x"ff760e79";
		wait for Clk_period;
		Addr <=  "0001110010001";
		Trees_din <= x"000cd30c";
		wait for Clk_period;
		Addr <=  "0001110010010";
		Trees_din <= x"000c8b08";
		wait for Clk_period;
		Addr <=  "0001110010011";
		Trees_din <= x"07fb0a04";
		wait for Clk_period;
		Addr <=  "0001110010100";
		Trees_din <= x"ffde0e79";
		wait for Clk_period;
		Addr <=  "0001110010101";
		Trees_din <= x"006c0e79";
		wait for Clk_period;
		Addr <=  "0001110010110";
		Trees_din <= x"00ed0e79";
		wait for Clk_period;
		Addr <=  "0001110010111";
		Trees_din <= x"0408b408";
		wait for Clk_period;
		Addr <=  "0001110011000";
		Trees_din <= x"07fc7104";
		wait for Clk_period;
		Addr <=  "0001110011001";
		Trees_din <= x"ff780e79";
		wait for Clk_period;
		Addr <=  "0001110011010";
		Trees_din <= x"ffe30e79";
		wait for Clk_period;
		Addr <=  "0001110011011";
		Trees_din <= x"07f7cc04";
		wait for Clk_period;
		Addr <=  "0001110011100";
		Trees_din <= x"ffce0e79";
		wait for Clk_period;
		Addr <=  "0001110011101";
		Trees_din <= x"00670e79";
		wait for Clk_period;
		Addr <=  "0001110011110";
		Trees_din <= x"04ffbc2c";
		wait for Clk_period;
		Addr <=  "0001110011111";
		Trees_din <= x"010c6428";
		wait for Clk_period;
		Addr <=  "0001110100000";
		Trees_din <= x"0b006610";
		wait for Clk_period;
		Addr <=  "0001110100001";
		Trees_din <= x"05f5e008";
		wait for Clk_period;
		Addr <=  "0001110100010";
		Trees_din <= x"0e003504";
		wait for Clk_period;
		Addr <=  "0001110100011";
		Trees_din <= x"01760f3d";
		wait for Clk_period;
		Addr <=  "0001110100100";
		Trees_din <= x"ffb10f3d";
		wait for Clk_period;
		Addr <=  "0001110100101";
		Trees_din <= x"1afd9b04";
		wait for Clk_period;
		Addr <=  "0001110100110";
		Trees_din <= x"ff860f3d";
		wait for Clk_period;
		Addr <=  "0001110100111";
		Trees_din <= x"002a0f3d";
		wait for Clk_period;
		Addr <=  "0001110101000";
		Trees_din <= x"0f00020c";
		wait for Clk_period;
		Addr <=  "0001110101001";
		Trees_din <= x"10004208";
		wait for Clk_period;
		Addr <=  "0001110101010";
		Trees_din <= x"07012a04";
		wait for Clk_period;
		Addr <=  "0001110101011";
		Trees_din <= x"002e0f3d";
		wait for Clk_period;
		Addr <=  "0001110101100";
		Trees_din <= x"00d80f3d";
		wait for Clk_period;
		Addr <=  "0001110101101";
		Trees_din <= x"ff8f0f3d";
		wait for Clk_period;
		Addr <=  "0001110101110";
		Trees_din <= x"16004e08";
		wait for Clk_period;
		Addr <=  "0001110101111";
		Trees_din <= x"1100d204";
		wait for Clk_period;
		Addr <=  "0001110110000";
		Trees_din <= x"00470f3d";
		wait for Clk_period;
		Addr <=  "0001110110001";
		Trees_din <= x"ff990f3d";
		wait for Clk_period;
		Addr <=  "0001110110010";
		Trees_din <= x"ff6e0f3d";
		wait for Clk_period;
		Addr <=  "0001110110011";
		Trees_din <= x"ff6d0f3d";
		wait for Clk_period;
		Addr <=  "0001110110100";
		Trees_din <= x"03f50b10";
		wait for Clk_period;
		Addr <=  "0001110110101";
		Trees_din <= x"04ffdd04";
		wait for Clk_period;
		Addr <=  "0001110110110";
		Trees_din <= x"00580f3d";
		wait for Clk_period;
		Addr <=  "0001110110111";
		Trees_din <= x"04080d04";
		wait for Clk_period;
		Addr <=  "0001110111000";
		Trees_din <= x"ff760f3d";
		wait for Clk_period;
		Addr <=  "0001110111001";
		Trees_din <= x"07f76704";
		wait for Clk_period;
		Addr <=  "0001110111010";
		Trees_din <= x"00340f3d";
		wait for Clk_period;
		Addr <=  "0001110111011";
		Trees_din <= x"ffd50f3d";
		wait for Clk_period;
		Addr <=  "0001110111100";
		Trees_din <= x"010e3220";
		wait for Clk_period;
		Addr <=  "0001110111101";
		Trees_din <= x"0209bd10";
		wait for Clk_period;
		Addr <=  "0001110111110";
		Trees_din <= x"16005c08";
		wait for Clk_period;
		Addr <=  "0001110111111";
		Trees_din <= x"04063004";
		wait for Clk_period;
		Addr <=  "0001111000000";
		Trees_din <= x"ff970f3d";
		wait for Clk_period;
		Addr <=  "0001111000001";
		Trees_din <= x"005c0f3d";
		wait for Clk_period;
		Addr <=  "0001111000010";
		Trees_din <= x"0e002704";
		wait for Clk_period;
		Addr <=  "0001111000011";
		Trees_din <= x"00b70f3d";
		wait for Clk_period;
		Addr <=  "0001111000100";
		Trees_din <= x"002b0f3d";
		wait for Clk_period;
		Addr <=  "0001111000101";
		Trees_din <= x"01ffc908";
		wait for Clk_period;
		Addr <=  "0001111000110";
		Trees_din <= x"10004504";
		wait for Clk_period;
		Addr <=  "0001111000111";
		Trees_din <= x"00990f3d";
		wait for Clk_period;
		Addr <=  "0001111001000";
		Trees_din <= x"ffe30f3d";
		wait for Clk_period;
		Addr <=  "0001111001001";
		Trees_din <= x"04057d04";
		wait for Clk_period;
		Addr <=  "0001111001010";
		Trees_din <= x"ff7a0f3d";
		wait for Clk_period;
		Addr <=  "0001111001011";
		Trees_din <= x"fff50f3d";
		wait for Clk_period;
		Addr <=  "0001111001100";
		Trees_din <= x"0c00bb04";
		wait for Clk_period;
		Addr <=  "0001111001101";
		Trees_din <= x"ff7b0f3d";
		wait for Clk_period;
		Addr <=  "0001111001110";
		Trees_din <= x"00330f3d";
		wait for Clk_period;
		Addr <=  "0001111001111";
		Trees_din <= x"04ff7c28";
		wait for Clk_period;
		Addr <=  "0001111010000";
		Trees_din <= x"0b006614";
		wait for Clk_period;
		Addr <=  "0001111010001";
		Trees_din <= x"0f001508";
		wait for Clk_period;
		Addr <=  "0001111010010";
		Trees_din <= x"13040004";
		wait for Clk_period;
		Addr <=  "0001111010011";
		Trees_din <= x"ff7b1021";
		wait for Clk_period;
		Addr <=  "0001111010100";
		Trees_din <= x"00211021";
		wait for Clk_period;
		Addr <=  "0001111010101";
		Trees_din <= x"0f002404";
		wait for Clk_period;
		Addr <=  "0001111010110";
		Trees_din <= x"01341021";
		wait for Clk_period;
		Addr <=  "0001111010111";
		Trees_din <= x"19000a04";
		wait for Clk_period;
		Addr <=  "0001111011000";
		Trees_din <= x"ffa21021";
		wait for Clk_period;
		Addr <=  "0001111011001";
		Trees_din <= x"001f1021";
		wait for Clk_period;
		Addr <=  "0001111011010";
		Trees_din <= x"0f000008";
		wait for Clk_period;
		Addr <=  "0001111011011";
		Trees_din <= x"11013704";
		wait for Clk_period;
		Addr <=  "0001111011100";
		Trees_din <= x"ff8f1021";
		wait for Clk_period;
		Addr <=  "0001111011101";
		Trees_din <= x"00c41021";
		wait for Clk_period;
		Addr <=  "0001111011110";
		Trees_din <= x"03fee004";
		wait for Clk_period;
		Addr <=  "0001111011111";
		Trees_din <= x"ff6b1021";
		wait for Clk_period;
		Addr <=  "0001111100000";
		Trees_din <= x"0c00c304";
		wait for Clk_period;
		Addr <=  "0001111100001";
		Trees_din <= x"ff8f1021";
		wait for Clk_period;
		Addr <=  "0001111100010";
		Trees_din <= x"003d1021";
		wait for Clk_period;
		Addr <=  "0001111100011";
		Trees_din <= x"0f00011c";
		wait for Clk_period;
		Addr <=  "0001111100100";
		Trees_din <= x"0c007c10";
		wait for Clk_period;
		Addr <=  "0001111100101";
		Trees_din <= x"0c006904";
		wait for Clk_period;
		Addr <=  "0001111100110";
		Trees_din <= x"ff9c1021";
		wait for Clk_period;
		Addr <=  "0001111100111";
		Trees_din <= x"06011908";
		wait for Clk_period;
		Addr <=  "0001111101000";
		Trees_din <= x"08004104";
		wait for Clk_period;
		Addr <=  "0001111101001";
		Trees_din <= x"002a1021";
		wait for Clk_period;
		Addr <=  "0001111101010";
		Trees_din <= x"00941021";
		wait for Clk_period;
		Addr <=  "0001111101011";
		Trees_din <= x"ffe81021";
		wait for Clk_period;
		Addr <=  "0001111101100";
		Trees_din <= x"0b009108";
		wait for Clk_period;
		Addr <=  "0001111101101";
		Trees_din <= x"1403fe04";
		wait for Clk_period;
		Addr <=  "0001111101110";
		Trees_din <= x"ffdd1021";
		wait for Clk_period;
		Addr <=  "0001111101111";
		Trees_din <= x"ff6e1021";
		wait for Clk_period;
		Addr <=  "0001111110000";
		Trees_din <= x"003a1021";
		wait for Clk_period;
		Addr <=  "0001111110001";
		Trees_din <= x"0f000414";
		wait for Clk_period;
		Addr <=  "0001111110010";
		Trees_din <= x"1403fe04";
		wait for Clk_period;
		Addr <=  "0001111110011";
		Trees_din <= x"ffab1021";
		wait for Clk_period;
		Addr <=  "0001111110100";
		Trees_din <= x"18002508";
		wait for Clk_period;
		Addr <=  "0001111110101";
		Trees_din <= x"0900ac04";
		wait for Clk_period;
		Addr <=  "0001111110110";
		Trees_din <= x"ffab1021";
		wait for Clk_period;
		Addr <=  "0001111110111";
		Trees_din <= x"00671021";
		wait for Clk_period;
		Addr <=  "0001111111000";
		Trees_din <= x"08003904";
		wait for Clk_period;
		Addr <=  "0001111111001";
		Trees_din <= x"00441021";
		wait for Clk_period;
		Addr <=  "0001111111010";
		Trees_din <= x"019b1021";
		wait for Clk_period;
		Addr <=  "0001111111011";
		Trees_din <= x"05f6af0c";
		wait for Clk_period;
		Addr <=  "0001111111100";
		Trees_din <= x"03fb4208";
		wait for Clk_period;
		Addr <=  "0001111111101";
		Trees_din <= x"000c2504";
		wait for Clk_period;
		Addr <=  "0001111111110";
		Trees_din <= x"ff901021";
		wait for Clk_period;
		Addr <=  "0001111111111";
		Trees_din <= x"fff91021";
		wait for Clk_period;
		Addr <=  "0010000000000";
		Trees_din <= x"00931021";
		wait for Clk_period;
		Addr <=  "0010000000001";
		Trees_din <= x"18004a08";
		wait for Clk_period;
		Addr <=  "0010000000010";
		Trees_din <= x"11001604";
		wait for Clk_period;
		Addr <=  "0010000000011";
		Trees_din <= x"00411021";
		wait for Clk_period;
		Addr <=  "0010000000100";
		Trees_din <= x"ff981021";
		wait for Clk_period;
		Addr <=  "0010000000101";
		Trees_din <= x"0c00af04";
		wait for Clk_period;
		Addr <=  "0010000000110";
		Trees_din <= x"00771021";
		wait for Clk_period;
		Addr <=  "0010000000111";
		Trees_din <= x"00031021";
		wait for Clk_period;
		Addr <=  "0010000001000";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0010000001001";
		Trees_din <= x"04ff7c24";
		wait for Clk_period;
		Addr <=  "0010000001010";
		Trees_din <= x"0d008d08";
		wait for Clk_period;
		Addr <=  "0010000001011";
		Trees_din <= x"0a003804";
		wait for Clk_period;
		Addr <=  "0010000001100";
		Trees_din <= x"00271111";
		wait for Clk_period;
		Addr <=  "0010000001101";
		Trees_din <= x"ff6d1111";
		wait for Clk_period;
		Addr <=  "0010000001110";
		Trees_din <= x"1403db08";
		wait for Clk_period;
		Addr <=  "0010000001111";
		Trees_din <= x"1c028704";
		wait for Clk_period;
		Addr <=  "0010000010000";
		Trees_din <= x"ff761111";
		wait for Clk_period;
		Addr <=  "0010000010001";
		Trees_din <= x"001d1111";
		wait for Clk_period;
		Addr <=  "0010000010010";
		Trees_din <= x"02054604";
		wait for Clk_period;
		Addr <=  "0010000010011";
		Trees_din <= x"ff851111";
		wait for Clk_period;
		Addr <=  "0010000010100";
		Trees_din <= x"0205e308";
		wait for Clk_period;
		Addr <=  "0010000010101";
		Trees_din <= x"04fbfc04";
		wait for Clk_period;
		Addr <=  "0010000010110";
		Trees_din <= x"01771111";
		wait for Clk_period;
		Addr <=  "0010000010111";
		Trees_din <= x"003c1111";
		wait for Clk_period;
		Addr <=  "0010000011000";
		Trees_din <= x"1800bc04";
		wait for Clk_period;
		Addr <=  "0010000011001";
		Trees_din <= x"ff991111";
		wait for Clk_period;
		Addr <=  "0010000011010";
		Trees_din <= x"00451111";
		wait for Clk_period;
		Addr <=  "0010000011011";
		Trees_din <= x"0900b824";
		wait for Clk_period;
		Addr <=  "0010000011100";
		Trees_din <= x"03f9c51c";
		wait for Clk_period;
		Addr <=  "0010000011101";
		Trees_din <= x"000ed010";
		wait for Clk_period;
		Addr <=  "0010000011110";
		Trees_din <= x"000de208";
		wait for Clk_period;
		Addr <=  "0010000011111";
		Trees_din <= x"1303a604";
		wait for Clk_period;
		Addr <=  "0010000100000";
		Trees_din <= x"ffdf1111";
		wait for Clk_period;
		Addr <=  "0010000100001";
		Trees_din <= x"00611111";
		wait for Clk_period;
		Addr <=  "0010000100010";
		Trees_din <= x"05f4da04";
		wait for Clk_period;
		Addr <=  "0010000100011";
		Trees_din <= x"ffed1111";
		wait for Clk_period;
		Addr <=  "0010000100100";
		Trees_din <= x"010d1111";
		wait for Clk_period;
		Addr <=  "0010000100101";
		Trees_din <= x"19002c08";
		wait for Clk_period;
		Addr <=  "0010000100110";
		Trees_din <= x"040a8404";
		wait for Clk_period;
		Addr <=  "0010000100111";
		Trees_din <= x"ff811111";
		wait for Clk_period;
		Addr <=  "0010000101000";
		Trees_din <= x"00161111";
		wait for Clk_period;
		Addr <=  "0010000101001";
		Trees_din <= x"005d1111";
		wait for Clk_period;
		Addr <=  "0010000101010";
		Trees_din <= x"0403e704";
		wait for Clk_period;
		Addr <=  "0010000101011";
		Trees_din <= x"ff851111";
		wait for Clk_period;
		Addr <=  "0010000101100";
		Trees_din <= x"000e1111";
		wait for Clk_period;
		Addr <=  "0010000101101";
		Trees_din <= x"0402ab14";
		wait for Clk_period;
		Addr <=  "0010000101110";
		Trees_din <= x"00123210";
		wait for Clk_period;
		Addr <=  "0010000101111";
		Trees_din <= x"1102cb08";
		wait for Clk_period;
		Addr <=  "0010000110000";
		Trees_din <= x"03fb4204";
		wait for Clk_period;
		Addr <=  "0010000110001";
		Trees_din <= x"ff781111";
		wait for Clk_period;
		Addr <=  "0010000110010";
		Trees_din <= x"00141111";
		wait for Clk_period;
		Addr <=  "0010000110011";
		Trees_din <= x"05f6dc04";
		wait for Clk_period;
		Addr <=  "0010000110100";
		Trees_din <= x"ffaf1111";
		wait for Clk_period;
		Addr <=  "0010000110101";
		Trees_din <= x"00911111";
		wait for Clk_period;
		Addr <=  "0010000110110";
		Trees_din <= x"00641111";
		wait for Clk_period;
		Addr <=  "0010000110111";
		Trees_din <= x"000d1b10";
		wait for Clk_period;
		Addr <=  "0010000111000";
		Trees_din <= x"02099108";
		wait for Clk_period;
		Addr <=  "0010000111001";
		Trees_din <= x"12007c04";
		wait for Clk_period;
		Addr <=  "0010000111010";
		Trees_din <= x"007c1111";
		wait for Clk_period;
		Addr <=  "0010000111011";
		Trees_din <= x"ffce1111";
		wait for Clk_period;
		Addr <=  "0010000111100";
		Trees_din <= x"10004104";
		wait for Clk_period;
		Addr <=  "0010000111101";
		Trees_din <= x"006d1111";
		wait for Clk_period;
		Addr <=  "0010000111110";
		Trees_din <= x"ff9d1111";
		wait for Clk_period;
		Addr <=  "0010000111111";
		Trees_din <= x"0408b404";
		wait for Clk_period;
		Addr <=  "0010001000000";
		Trees_din <= x"ff7f1111";
		wait for Clk_period;
		Addr <=  "0010001000001";
		Trees_din <= x"07f8d804";
		wait for Clk_period;
		Addr <=  "0010001000010";
		Trees_din <= x"ffd41111";
		wait for Clk_period;
		Addr <=  "0010001000011";
		Trees_din <= x"005c1111";
		wait for Clk_period;
		Addr <=  "0010001000100";
		Trees_din <= x"04ff7c24";
		wait for Clk_period;
		Addr <=  "0010001000101";
		Trees_din <= x"0b006614";
		wait for Clk_period;
		Addr <=  "0010001000110";
		Trees_din <= x"0f001508";
		wait for Clk_period;
		Addr <=  "0010001000111";
		Trees_din <= x"1600ab04";
		wait for Clk_period;
		Addr <=  "0010001001000";
		Trees_din <= x"ff8111f5";
		wait for Clk_period;
		Addr <=  "0010001001001";
		Trees_din <= x"002811f5";
		wait for Clk_period;
		Addr <=  "0010001001010";
		Trees_din <= x"0b006404";
		wait for Clk_period;
		Addr <=  "0010001001011";
		Trees_din <= x"ffa911f5";
		wait for Clk_period;
		Addr <=  "0010001001100";
		Trees_din <= x"0f002404";
		wait for Clk_period;
		Addr <=  "0010001001101";
		Trees_din <= x"011311f5";
		wait for Clk_period;
		Addr <=  "0010001001110";
		Trees_din <= x"001611f5";
		wait for Clk_period;
		Addr <=  "0010001001111";
		Trees_din <= x"03fee008";
		wait for Clk_period;
		Addr <=  "0010001010000";
		Trees_din <= x"01004904";
		wait for Clk_period;
		Addr <=  "0010001010001";
		Trees_din <= x"fff611f5";
		wait for Clk_period;
		Addr <=  "0010001010010";
		Trees_din <= x"ff6d11f5";
		wait for Clk_period;
		Addr <=  "0010001010011";
		Trees_din <= x"10004004";
		wait for Clk_period;
		Addr <=  "0010001010100";
		Trees_din <= x"008111f5";
		wait for Clk_period;
		Addr <=  "0010001010101";
		Trees_din <= x"ff9711f5";
		wait for Clk_period;
		Addr <=  "0010001010110";
		Trees_din <= x"0f00011c";
		wait for Clk_period;
		Addr <=  "0010001010111";
		Trees_din <= x"0c007c10";
		wait for Clk_period;
		Addr <=  "0010001011000";
		Trees_din <= x"0c006904";
		wait for Clk_period;
		Addr <=  "0010001011001";
		Trees_din <= x"ffa311f5";
		wait for Clk_period;
		Addr <=  "0010001011010";
		Trees_din <= x"10005404";
		wait for Clk_period;
		Addr <=  "0010001011011";
		Trees_din <= x"000511f5";
		wait for Clk_period;
		Addr <=  "0010001011100";
		Trees_din <= x"0a004504";
		wait for Clk_period;
		Addr <=  "0010001011101";
		Trees_din <= x"009111f5";
		wait for Clk_period;
		Addr <=  "0010001011110";
		Trees_din <= x"002011f5";
		wait for Clk_period;
		Addr <=  "0010001011111";
		Trees_din <= x"08003004";
		wait for Clk_period;
		Addr <=  "0010001100000";
		Trees_din <= x"003111f5";
		wait for Clk_period;
		Addr <=  "0010001100001";
		Trees_din <= x"01fed304";
		wait for Clk_period;
		Addr <=  "0010001100010";
		Trees_din <= x"ffe611f5";
		wait for Clk_period;
		Addr <=  "0010001100011";
		Trees_din <= x"ff7111f5";
		wait for Clk_period;
		Addr <=  "0010001100100";
		Trees_din <= x"0f000414";
		wait for Clk_period;
		Addr <=  "0010001100101";
		Trees_din <= x"10005010";
		wait for Clk_period;
		Addr <=  "0010001100110";
		Trees_din <= x"0900b508";
		wait for Clk_period;
		Addr <=  "0010001100111";
		Trees_din <= x"0900ad04";
		wait for Clk_period;
		Addr <=  "0010001101000";
		Trees_din <= x"005611f5";
		wait for Clk_period;
		Addr <=  "0010001101001";
		Trees_din <= x"00fc11f5";
		wait for Clk_period;
		Addr <=  "0010001101010";
		Trees_din <= x"0403d204";
		wait for Clk_period;
		Addr <=  "0010001101011";
		Trees_din <= x"ffaa11f5";
		wait for Clk_period;
		Addr <=  "0010001101100";
		Trees_din <= x"006611f5";
		wait for Clk_period;
		Addr <=  "0010001101101";
		Trees_din <= x"ffc811f5";
		wait for Clk_period;
		Addr <=  "0010001101110";
		Trees_din <= x"010b6e10";
		wait for Clk_period;
		Addr <=  "0010001101111";
		Trees_din <= x"0900ec08";
		wait for Clk_period;
		Addr <=  "0010001110000";
		Trees_din <= x"03f50b04";
		wait for Clk_period;
		Addr <=  "0010001110001";
		Trees_din <= x"ff9e11f5";
		wait for Clk_period;
		Addr <=  "0010001110010";
		Trees_din <= x"003211f5";
		wait for Clk_period;
		Addr <=  "0010001110011";
		Trees_din <= x"03f52504";
		wait for Clk_period;
		Addr <=  "0010001110100";
		Trees_din <= x"003a11f5";
		wait for Clk_period;
		Addr <=  "0010001110101";
		Trees_din <= x"ff7a11f5";
		wait for Clk_period;
		Addr <=  "0010001110110";
		Trees_din <= x"1c028708";
		wait for Clk_period;
		Addr <=  "0010001110111";
		Trees_din <= x"04032304";
		wait for Clk_period;
		Addr <=  "0010001111000";
		Trees_din <= x"ff7411f5";
		wait for Clk_period;
		Addr <=  "0010001111001";
		Trees_din <= x"fff511f5";
		wait for Clk_period;
		Addr <=  "0010001111010";
		Trees_din <= x"0e003204";
		wait for Clk_period;
		Addr <=  "0010001111011";
		Trees_din <= x"002211f5";
		wait for Clk_period;
		Addr <=  "0010001111100";
		Trees_din <= x"008c11f5";
		wait for Clk_period;
		Addr <=  "0010001111101";
		Trees_din <= x"04ffbc28";
		wait for Clk_period;
		Addr <=  "0010001111110";
		Trees_din <= x"010c6424";
		wait for Clk_period;
		Addr <=  "0010001111111";
		Trees_din <= x"0b00660c";
		wait for Clk_period;
		Addr <=  "0010010000000";
		Trees_din <= x"05f6cc08";
		wait for Clk_period;
		Addr <=  "0010010000001";
		Trees_din <= x"0f001404";
		wait for Clk_period;
		Addr <=  "0010010000010";
		Trees_din <= x"fff81311";
		wait for Clk_period;
		Addr <=  "0010010000011";
		Trees_din <= x"00d71311";
		wait for Clk_period;
		Addr <=  "0010010000100";
		Trees_din <= x"ff971311";
		wait for Clk_period;
		Addr <=  "0010010000101";
		Trees_din <= x"0f00020c";
		wait for Clk_period;
		Addr <=  "0010010000110";
		Trees_din <= x"10004208";
		wait for Clk_period;
		Addr <=  "0010010000111";
		Trees_din <= x"1303c304";
		wait for Clk_period;
		Addr <=  "0010010001000";
		Trees_din <= x"00ba1311";
		wait for Clk_period;
		Addr <=  "0010010001001";
		Trees_din <= x"00181311";
		wait for Clk_period;
		Addr <=  "0010010001010";
		Trees_din <= x"ffa01311";
		wait for Clk_period;
		Addr <=  "0010010001011";
		Trees_din <= x"16004e08";
		wait for Clk_period;
		Addr <=  "0010010001100";
		Trees_din <= x"0a004104";
		wait for Clk_period;
		Addr <=  "0010010001101";
		Trees_din <= x"ffae1311";
		wait for Clk_period;
		Addr <=  "0010010001110";
		Trees_din <= x"00421311";
		wait for Clk_period;
		Addr <=  "0010010001111";
		Trees_din <= x"ff751311";
		wait for Clk_period;
		Addr <=  "0010010010000";
		Trees_din <= x"ff731311";
		wait for Clk_period;
		Addr <=  "0010010010001";
		Trees_din <= x"08004138";
		wait for Clk_period;
		Addr <=  "0010010010010";
		Trees_din <= x"11015b18";
		wait for Clk_period;
		Addr <=  "0010010010011";
		Trees_din <= x"0d00000c";
		wait for Clk_period;
		Addr <=  "0010010010100";
		Trees_din <= x"0e002b08";
		wait for Clk_period;
		Addr <=  "0010010010101";
		Trees_din <= x"0e002104";
		wait for Clk_period;
		Addr <=  "0010010010110";
		Trees_din <= x"00001311";
		wait for Clk_period;
		Addr <=  "0010010010111";
		Trees_din <= x"00761311";
		wait for Clk_period;
		Addr <=  "0010010011000";
		Trees_din <= x"ff9e1311";
		wait for Clk_period;
		Addr <=  "0010010011001";
		Trees_din <= x"0403e704";
		wait for Clk_period;
		Addr <=  "0010010011010";
		Trees_din <= x"ff711311";
		wait for Clk_period;
		Addr <=  "0010010011011";
		Trees_din <= x"17f70f04";
		wait for Clk_period;
		Addr <=  "0010010011100";
		Trees_din <= x"00551311";
		wait for Clk_period;
		Addr <=  "0010010011101";
		Trees_din <= x"ffc01311";
		wait for Clk_period;
		Addr <=  "0010010011110";
		Trees_din <= x"16006d10";
		wait for Clk_period;
		Addr <=  "0010010011111";
		Trees_din <= x"0e002708";
		wait for Clk_period;
		Addr <=  "0010010100000";
		Trees_din <= x"0b007d04";
		wait for Clk_period;
		Addr <=  "0010010100001";
		Trees_din <= x"00ae1311";
		wait for Clk_period;
		Addr <=  "0010010100010";
		Trees_din <= x"ffd61311";
		wait for Clk_period;
		Addr <=  "0010010100011";
		Trees_din <= x"05f7fb04";
		wait for Clk_period;
		Addr <=  "0010010100100";
		Trees_din <= x"ff831311";
		wait for Clk_period;
		Addr <=  "0010010100101";
		Trees_din <= x"00031311";
		wait for Clk_period;
		Addr <=  "0010010100110";
		Trees_din <= x"08003c08";
		wait for Clk_period;
		Addr <=  "0010010100111";
		Trees_din <= x"05f75104";
		wait for Clk_period;
		Addr <=  "0010010101000";
		Trees_din <= x"00db1311";
		wait for Clk_period;
		Addr <=  "0010010101001";
		Trees_din <= x"00161311";
		wait for Clk_period;
		Addr <=  "0010010101010";
		Trees_din <= x"01079704";
		wait for Clk_period;
		Addr <=  "0010010101011";
		Trees_din <= x"00431311";
		wait for Clk_period;
		Addr <=  "0010010101100";
		Trees_din <= x"ffaf1311";
		wait for Clk_period;
		Addr <=  "0010010101101";
		Trees_din <= x"0800431c";
		wait for Clk_period;
		Addr <=  "0010010101110";
		Trees_din <= x"0d00b710";
		wait for Clk_period;
		Addr <=  "0010010101111";
		Trees_din <= x"1e026508";
		wait for Clk_period;
		Addr <=  "0010010110000";
		Trees_din <= x"04033e04";
		wait for Clk_period;
		Addr <=  "0010010110001";
		Trees_din <= x"ffad1311";
		wait for Clk_period;
		Addr <=  "0010010110010";
		Trees_din <= x"00761311";
		wait for Clk_period;
		Addr <=  "0010010110011";
		Trees_din <= x"10004104";
		wait for Clk_period;
		Addr <=  "0010010110100";
		Trees_din <= x"01601311";
		wait for Clk_period;
		Addr <=  "0010010110101";
		Trees_din <= x"005e1311";
		wait for Clk_period;
		Addr <=  "0010010110110";
		Trees_din <= x"1e027b04";
		wait for Clk_period;
		Addr <=  "0010010110111";
		Trees_din <= x"ffa01311";
		wait for Clk_period;
		Addr <=  "0010010111000";
		Trees_din <= x"05f66804";
		wait for Clk_period;
		Addr <=  "0010010111001";
		Trees_din <= x"00041311";
		wait for Clk_period;
		Addr <=  "0010010111010";
		Trees_din <= x"00851311";
		wait for Clk_period;
		Addr <=  "0010010111011";
		Trees_din <= x"03f9c510";
		wait for Clk_period;
		Addr <=  "0010010111100";
		Trees_din <= x"1303cb08";
		wait for Clk_period;
		Addr <=  "0010010111101";
		Trees_din <= x"0d01f704";
		wait for Clk_period;
		Addr <=  "0010010111110";
		Trees_din <= x"ffb21311";
		wait for Clk_period;
		Addr <=  "0010010111111";
		Trees_din <= x"00251311";
		wait for Clk_period;
		Addr <=  "0010011000000";
		Trees_din <= x"10004c04";
		wait for Clk_period;
		Addr <=  "0010011000001";
		Trees_din <= x"00751311";
		wait for Clk_period;
		Addr <=  "0010011000010";
		Trees_din <= x"ffe81311";
		wait for Clk_period;
		Addr <=  "0010011000011";
		Trees_din <= x"ff7b1311";
		wait for Clk_period;
		Addr <=  "0010011000100";
		Trees_din <= x"04ff7c20";
		wait for Clk_period;
		Addr <=  "0010011000101";
		Trees_din <= x"02054608";
		wait for Clk_period;
		Addr <=  "0010011000110";
		Trees_din <= x"1b028704";
		wait for Clk_period;
		Addr <=  "0010011000111";
		Trees_din <= x"ff7213d5";
		wait for Clk_period;
		Addr <=  "0010011001000";
		Trees_din <= x"000e13d5";
		wait for Clk_period;
		Addr <=  "0010011001001";
		Trees_din <= x"0205e30c";
		wait for Clk_period;
		Addr <=  "0010011001010";
		Trees_din <= x"07ffe904";
		wait for Clk_period;
		Addr <=  "0010011001011";
		Trees_din <= x"ffaa13d5";
		wait for Clk_period;
		Addr <=  "0010011001100";
		Trees_din <= x"04fbfc04";
		wait for Clk_period;
		Addr <=  "0010011001101";
		Trees_din <= x"00f113d5";
		wait for Clk_period;
		Addr <=  "0010011001110";
		Trees_din <= x"003313d5";
		wait for Clk_period;
		Addr <=  "0010011001111";
		Trees_din <= x"0b006408";
		wait for Clk_period;
		Addr <=  "0010011010000";
		Trees_din <= x"010b2804";
		wait for Clk_period;
		Addr <=  "0010011010001";
		Trees_din <= x"ffac13d5";
		wait for Clk_period;
		Addr <=  "0010011010010";
		Trees_din <= x"007713d5";
		wait for Clk_period;
		Addr <=  "0010011010011";
		Trees_din <= x"ff7713d5";
		wait for Clk_period;
		Addr <=  "0010011010100";
		Trees_din <= x"04057d2c";
		wait for Clk_period;
		Addr <=  "0010011010101";
		Trees_din <= x"06015b14";
		wait for Clk_period;
		Addr <=  "0010011010110";
		Trees_din <= x"16005c04";
		wait for Clk_period;
		Addr <=  "0010011010111";
		Trees_din <= x"ff7f13d5";
		wait for Clk_period;
		Addr <=  "0010011011000";
		Trees_din <= x"0c009e08";
		wait for Clk_period;
		Addr <=  "0010011011001";
		Trees_din <= x"06010c04";
		wait for Clk_period;
		Addr <=  "0010011011010";
		Trees_din <= x"ffc413d5";
		wait for Clk_period;
		Addr <=  "0010011011011";
		Trees_din <= x"007f13d5";
		wait for Clk_period;
		Addr <=  "0010011011100";
		Trees_din <= x"02083304";
		wait for Clk_period;
		Addr <=  "0010011011101";
		Trees_din <= x"005e13d5";
		wait for Clk_period;
		Addr <=  "0010011011110";
		Trees_din <= x"ffc113d5";
		wait for Clk_period;
		Addr <=  "0010011011111";
		Trees_din <= x"15003d10";
		wait for Clk_period;
		Addr <=  "0010011100000";
		Trees_din <= x"07fd5f08";
		wait for Clk_period;
		Addr <=  "0010011100001";
		Trees_din <= x"0403e704";
		wait for Clk_period;
		Addr <=  "0010011100010";
		Trees_din <= x"ff8513d5";
		wait for Clk_period;
		Addr <=  "0010011100011";
		Trees_din <= x"001f13d5";
		wait for Clk_period;
		Addr <=  "0010011100100";
		Trees_din <= x"1afbd904";
		wait for Clk_period;
		Addr <=  "0010011100101";
		Trees_din <= x"008913d5";
		wait for Clk_period;
		Addr <=  "0010011100110";
		Trees_din <= x"000013d5";
		wait for Clk_period;
		Addr <=  "0010011100111";
		Trees_din <= x"010d4c04";
		wait for Clk_period;
		Addr <=  "0010011101000";
		Trees_din <= x"ff6c13d5";
		wait for Clk_period;
		Addr <=  "0010011101001";
		Trees_din <= x"000113d5";
		wait for Clk_period;
		Addr <=  "0010011101010";
		Trees_din <= x"0109ed14";
		wait for Clk_period;
		Addr <=  "0010011101011";
		Trees_din <= x"020d790c";
		wait for Clk_period;
		Addr <=  "0010011101100";
		Trees_din <= x"1102b608";
		wait for Clk_period;
		Addr <=  "0010011101101";
		Trees_din <= x"18001704";
		wait for Clk_period;
		Addr <=  "0010011101110";
		Trees_din <= x"fff213d5";
		wait for Clk_period;
		Addr <=  "0010011101111";
		Trees_din <= x"008113d5";
		wait for Clk_period;
		Addr <=  "0010011110000";
		Trees_din <= x"ffd613d5";
		wait for Clk_period;
		Addr <=  "0010011110001";
		Trees_din <= x"01fdba04";
		wait for Clk_period;
		Addr <=  "0010011110010";
		Trees_din <= x"001513d5";
		wait for Clk_period;
		Addr <=  "0010011110011";
		Trees_din <= x"ffa913d5";
		wait for Clk_period;
		Addr <=  "0010011110100";
		Trees_din <= x"ff9b13d5";
		wait for Clk_period;
		Addr <=  "0010011110101";
		Trees_din <= x"04001728";
		wait for Clk_period;
		Addr <=  "0010011110110";
		Trees_din <= x"06ff080c";
		wait for Clk_period;
		Addr <=  "0010011110111";
		Trees_din <= x"1102d808";
		wait for Clk_period;
		Addr <=  "0010011111000";
		Trees_din <= x"1e028704";
		wait for Clk_period;
		Addr <=  "0010011111001";
		Trees_din <= x"ff731479";
		wait for Clk_period;
		Addr <=  "0010011111010";
		Trees_din <= x"fffb1479";
		wait for Clk_period;
		Addr <=  "0010011111011";
		Trees_din <= x"00261479";
		wait for Clk_period;
		Addr <=  "0010011111100";
		Trees_din <= x"06ff3f04";
		wait for Clk_period;
		Addr <=  "0010011111101";
		Trees_din <= x"00761479";
		wait for Clk_period;
		Addr <=  "0010011111110";
		Trees_din <= x"0b00690c";
		wait for Clk_period;
		Addr <=  "0010011111111";
		Trees_din <= x"05f6cc08";
		wait for Clk_period;
		Addr <=  "0010100000000";
		Trees_din <= x"0205e304";
		wait for Clk_period;
		Addr <=  "0010100000001";
		Trees_din <= x"00881479";
		wait for Clk_period;
		Addr <=  "0010100000010";
		Trees_din <= x"ffe51479";
		wait for Clk_period;
		Addr <=  "0010100000011";
		Trees_din <= x"ff9e1479";
		wait for Clk_period;
		Addr <=  "0010100000100";
		Trees_din <= x"0b008b04";
		wait for Clk_period;
		Addr <=  "0010100000101";
		Trees_din <= x"ff791479";
		wait for Clk_period;
		Addr <=  "0010100000110";
		Trees_din <= x"17f78504";
		wait for Clk_period;
		Addr <=  "0010100000111";
		Trees_din <= x"00651479";
		wait for Clk_period;
		Addr <=  "0010100001000";
		Trees_din <= x"ffaa1479";
		wait for Clk_period;
		Addr <=  "0010100001001";
		Trees_din <= x"03f50b08";
		wait for Clk_period;
		Addr <=  "0010100001010";
		Trees_din <= x"00098404";
		wait for Clk_period;
		Addr <=  "0010100001011";
		Trees_din <= x"00241479";
		wait for Clk_period;
		Addr <=  "0010100001100";
		Trees_din <= x"ff8d1479";
		wait for Clk_period;
		Addr <=  "0010100001101";
		Trees_din <= x"13018a04";
		wait for Clk_period;
		Addr <=  "0010100001110";
		Trees_din <= x"ff931479";
		wait for Clk_period;
		Addr <=  "0010100001111";
		Trees_din <= x"03f5e510";
		wait for Clk_period;
		Addr <=  "0010100010000";
		Trees_din <= x"0d006d08";
		wait for Clk_period;
		Addr <=  "0010100010001";
		Trees_din <= x"0603ba04";
		wait for Clk_period;
		Addr <=  "0010100010010";
		Trees_din <= x"ffc91479";
		wait for Clk_period;
		Addr <=  "0010100010011";
		Trees_din <= x"003c1479";
		wait for Clk_period;
		Addr <=  "0010100010100";
		Trees_din <= x"07f9b904";
		wait for Clk_period;
		Addr <=  "0010100010101";
		Trees_din <= x"fff61479";
		wait for Clk_period;
		Addr <=  "0010100010110";
		Trees_din <= x"00dc1479";
		wait for Clk_period;
		Addr <=  "0010100010111";
		Trees_din <= x"13022b08";
		wait for Clk_period;
		Addr <=  "0010100011000";
		Trees_din <= x"05f56804";
		wait for Clk_period;
		Addr <=  "0010100011001";
		Trees_din <= x"ffd11479";
		wait for Clk_period;
		Addr <=  "0010100011010";
		Trees_din <= x"008f1479";
		wait for Clk_period;
		Addr <=  "0010100011011";
		Trees_din <= x"11028f04";
		wait for Clk_period;
		Addr <=  "0010100011100";
		Trees_din <= x"000b1479";
		wait for Clk_period;
		Addr <=  "0010100011101";
		Trees_din <= x"ff921479";
		wait for Clk_period;
		Addr <=  "0010100011110";
		Trees_din <= x"04032338";
		wait for Clk_period;
		Addr <=  "0010100011111";
		Trees_din <= x"0c00950c";
		wait for Clk_period;
		Addr <=  "0010100100000";
		Trees_din <= x"14040004";
		wait for Clk_period;
		Addr <=  "0010100100001";
		Trees_din <= x"ff761575";
		wait for Clk_period;
		Addr <=  "0010100100010";
		Trees_din <= x"0a004504";
		wait for Clk_period;
		Addr <=  "0010100100011";
		Trees_din <= x"00441575";
		wait for Clk_period;
		Addr <=  "0010100100100";
		Trees_din <= x"ffa71575";
		wait for Clk_period;
		Addr <=  "0010100100101";
		Trees_din <= x"0d00000c";
		wait for Clk_period;
		Addr <=  "0010100100110";
		Trees_din <= x"1afbf808";
		wait for Clk_period;
		Addr <=  "0010100100111";
		Trees_din <= x"08003f04";
		wait for Clk_period;
		Addr <=  "0010100101000";
		Trees_din <= x"00261575";
		wait for Clk_period;
		Addr <=  "0010100101001";
		Trees_din <= x"00c81575";
		wait for Clk_period;
		Addr <=  "0010100101010";
		Trees_din <= x"ffeb1575";
		wait for Clk_period;
		Addr <=  "0010100101011";
		Trees_din <= x"0e003210";
		wait for Clk_period;
		Addr <=  "0010100101100";
		Trees_din <= x"16006d08";
		wait for Clk_period;
		Addr <=  "0010100101101";
		Trees_din <= x"16006004";
		wait for Clk_period;
		Addr <=  "0010100101110";
		Trees_din <= x"ffd91575";
		wait for Clk_period;
		Addr <=  "0010100101111";
		Trees_din <= x"ff731575";
		wait for Clk_period;
		Addr <=  "0010100110000";
		Trees_din <= x"16006d04";
		wait for Clk_period;
		Addr <=  "0010100110001";
		Trees_din <= x"00b51575";
		wait for Clk_period;
		Addr <=  "0010100110010";
		Trees_din <= x"ffd91575";
		wait for Clk_period;
		Addr <=  "0010100110011";
		Trees_din <= x"10004208";
		wait for Clk_period;
		Addr <=  "0010100110100";
		Trees_din <= x"11011e04";
		wait for Clk_period;
		Addr <=  "0010100110101";
		Trees_din <= x"001d1575";
		wait for Clk_period;
		Addr <=  "0010100110110";
		Trees_din <= x"00c81575";
		wait for Clk_period;
		Addr <=  "0010100110111";
		Trees_din <= x"0b006904";
		wait for Clk_period;
		Addr <=  "0010100111000";
		Trees_din <= x"00331575";
		wait for Clk_period;
		Addr <=  "0010100111001";
		Trees_din <= x"ffaa1575";
		wait for Clk_period;
		Addr <=  "0010100111010";
		Trees_din <= x"10004828";
		wait for Clk_period;
		Addr <=  "0010100111011";
		Trees_din <= x"0d008510";
		wait for Clk_period;
		Addr <=  "0010100111100";
		Trees_din <= x"040a840c";
		wait for Clk_period;
		Addr <=  "0010100111101";
		Trees_din <= x"0e001f04";
		wait for Clk_period;
		Addr <=  "0010100111110";
		Trees_din <= x"00221575";
		wait for Clk_period;
		Addr <=  "0010100111111";
		Trees_din <= x"07fc0d04";
		wait for Clk_period;
		Addr <=  "0010101000000";
		Trees_din <= x"ff6f1575";
		wait for Clk_period;
		Addr <=  "0010101000001";
		Trees_din <= x"fff21575";
		wait for Clk_period;
		Addr <=  "0010101000010";
		Trees_din <= x"00441575";
		wait for Clk_period;
		Addr <=  "0010101000011";
		Trees_din <= x"03f8310c";
		wait for Clk_period;
		Addr <=  "0010101000100";
		Trees_din <= x"06feca04";
		wait for Clk_period;
		Addr <=  "0010101000101";
		Trees_din <= x"003f1575";
		wait for Clk_period;
		Addr <=  "0010101000110";
		Trees_din <= x"11020e04";
		wait for Clk_period;
		Addr <=  "0010101000111";
		Trees_din <= x"ff9a1575";
		wait for Clk_period;
		Addr <=  "0010101001000";
		Trees_din <= x"fff11575";
		wait for Clk_period;
		Addr <=  "0010101001001";
		Trees_din <= x"08004208";
		wait for Clk_period;
		Addr <=  "0010101001010";
		Trees_din <= x"0b007204";
		wait for Clk_period;
		Addr <=  "0010101001011";
		Trees_din <= x"00351575";
		wait for Clk_period;
		Addr <=  "0010101001100";
		Trees_din <= x"00a51575";
		wait for Clk_period;
		Addr <=  "0010101001101";
		Trees_din <= x"ffec1575";
		wait for Clk_period;
		Addr <=  "0010101001110";
		Trees_din <= x"020b0318";
		wait for Clk_period;
		Addr <=  "0010101001111";
		Trees_din <= x"000e8010";
		wait for Clk_period;
		Addr <=  "0010101010000";
		Trees_din <= x"05f4e008";
		wait for Clk_period;
		Addr <=  "0010101010001";
		Trees_din <= x"1303d604";
		wait for Clk_period;
		Addr <=  "0010101010010";
		Trees_din <= x"ffcf1575";
		wait for Clk_period;
		Addr <=  "0010101010011";
		Trees_din <= x"00321575";
		wait for Clk_period;
		Addr <=  "0010101010100";
		Trees_din <= x"03f76604";
		wait for Clk_period;
		Addr <=  "0010101010101";
		Trees_din <= x"003b1575";
		wait for Clk_period;
		Addr <=  "0010101010110";
		Trees_din <= x"009d1575";
		wait for Clk_period;
		Addr <=  "0010101010111";
		Trees_din <= x"07f88604";
		wait for Clk_period;
		Addr <=  "0010101011000";
		Trees_din <= x"ffa61575";
		wait for Clk_period;
		Addr <=  "0010101011001";
		Trees_din <= x"00401575";
		wait for Clk_period;
		Addr <=  "0010101011010";
		Trees_din <= x"04098204";
		wait for Clk_period;
		Addr <=  "0010101011011";
		Trees_din <= x"ff951575";
		wait for Clk_period;
		Addr <=  "0010101011100";
		Trees_din <= x"001b1575";
		wait for Clk_period;
		Addr <=  "0010101011101";
		Trees_din <= x"010ce344";
		wait for Clk_period;
		Addr <=  "0010101011110";
		Trees_din <= x"06034b24";
		wait for Clk_period;
		Addr <=  "0010101011111";
		Trees_din <= x"05faad18";
		wait for Clk_period;
		Addr <=  "0010101100000";
		Trees_din <= x"15003008";
		wait for Clk_period;
		Addr <=  "0010101100001";
		Trees_din <= x"07f8b704";
		wait for Clk_period;
		Addr <=  "0010101100010";
		Trees_din <= x"fff51629";
		wait for Clk_period;
		Addr <=  "0010101100011";
		Trees_din <= x"ff8e1629";
		wait for Clk_period;
		Addr <=  "0010101100100";
		Trees_din <= x"02076e08";
		wait for Clk_period;
		Addr <=  "0010101100101";
		Trees_din <= x"08004a04";
		wait for Clk_period;
		Addr <=  "0010101100110";
		Trees_din <= x"005b1629";
		wait for Clk_period;
		Addr <=  "0010101100111";
		Trees_din <= x"ff961629";
		wait for Clk_period;
		Addr <=  "0010101101000";
		Trees_din <= x"04009f04";
		wait for Clk_period;
		Addr <=  "0010101101001";
		Trees_din <= x"ff891629";
		wait for Clk_period;
		Addr <=  "0010101101010";
		Trees_din <= x"001b1629";
		wait for Clk_period;
		Addr <=  "0010101101011";
		Trees_din <= x"0403fc04";
		wait for Clk_period;
		Addr <=  "0010101101100";
		Trees_din <= x"ff861629";
		wait for Clk_period;
		Addr <=  "0010101101101";
		Trees_din <= x"07fb6804";
		wait for Clk_period;
		Addr <=  "0010101101110";
		Trees_din <= x"ffc71629";
		wait for Clk_period;
		Addr <=  "0010101101111";
		Trees_din <= x"00391629";
		wait for Clk_period;
		Addr <=  "0010101110000";
		Trees_din <= x"01ffc910";
		wait for Clk_period;
		Addr <=  "0010101110001";
		Trees_din <= x"10004208";
		wait for Clk_period;
		Addr <=  "0010101110010";
		Trees_din <= x"0c00b604";
		wait for Clk_period;
		Addr <=  "0010101110011";
		Trees_din <= x"00871629";
		wait for Clk_period;
		Addr <=  "0010101110100";
		Trees_din <= x"ffec1629";
		wait for Clk_period;
		Addr <=  "0010101110101";
		Trees_din <= x"15004404";
		wait for Clk_period;
		Addr <=  "0010101110110";
		Trees_din <= x"ffab1629";
		wait for Clk_period;
		Addr <=  "0010101110111";
		Trees_din <= x"00021629";
		wait for Clk_period;
		Addr <=  "0010101111000";
		Trees_din <= x"07f6b404";
		wait for Clk_period;
		Addr <=  "0010101111001";
		Trees_din <= x"00361629";
		wait for Clk_period;
		Addr <=  "0010101111010";
		Trees_din <= x"10003d04";
		wait for Clk_period;
		Addr <=  "0010101111011";
		Trees_din <= x"ffdd1629";
		wait for Clk_period;
		Addr <=  "0010101111100";
		Trees_din <= x"1b028504";
		wait for Clk_period;
		Addr <=  "0010101111101";
		Trees_din <= x"ff761629";
		wait for Clk_period;
		Addr <=  "0010101111110";
		Trees_din <= x"ffd91629";
		wait for Clk_period;
		Addr <=  "0010101111111";
		Trees_din <= x"1c028710";
		wait for Clk_period;
		Addr <=  "0010110000000";
		Trees_din <= x"06034b0c";
		wait for Clk_period;
		Addr <=  "0010110000001";
		Trees_din <= x"0c00bd04";
		wait for Clk_period;
		Addr <=  "0010110000010";
		Trees_din <= x"ff711629";
		wait for Clk_period;
		Addr <=  "0010110000011";
		Trees_din <= x"0e003204";
		wait for Clk_period;
		Addr <=  "0010110000100";
		Trees_din <= x"ff921629";
		wait for Clk_period;
		Addr <=  "0010110000101";
		Trees_din <= x"005d1629";
		wait for Clk_period;
		Addr <=  "0010110000110";
		Trees_din <= x"00321629";
		wait for Clk_period;
		Addr <=  "0010110000111";
		Trees_din <= x"0d001504";
		wait for Clk_period;
		Addr <=  "0010110001000";
		Trees_din <= x"00761629";
		wait for Clk_period;
		Addr <=  "0010110001001";
		Trees_din <= x"001d1629";
		wait for Clk_period;
		Addr <=  "0010110001010";
		Trees_din <= x"04032338";
		wait for Clk_period;
		Addr <=  "0010110001011";
		Trees_din <= x"0c00950c";
		wait for Clk_period;
		Addr <=  "0010110001100";
		Trees_din <= x"14040004";
		wait for Clk_period;
		Addr <=  "0010110001101";
		Trees_din <= x"ff79170d";
		wait for Clk_period;
		Addr <=  "0010110001110";
		Trees_din <= x"0a004504";
		wait for Clk_period;
		Addr <=  "0010110001111";
		Trees_din <= x"0037170d";
		wait for Clk_period;
		Addr <=  "0010110010000";
		Trees_din <= x"ffae170d";
		wait for Clk_period;
		Addr <=  "0010110010001";
		Trees_din <= x"0d00000c";
		wait for Clk_period;
		Addr <=  "0010110010010";
		Trees_din <= x"1c027804";
		wait for Clk_period;
		Addr <=  "0010110010011";
		Trees_din <= x"fff5170d";
		wait for Clk_period;
		Addr <=  "0010110010100";
		Trees_din <= x"17f86104";
		wait for Clk_period;
		Addr <=  "0010110010101";
		Trees_din <= x"00b5170d";
		wait for Clk_period;
		Addr <=  "0010110010110";
		Trees_din <= x"002a170d";
		wait for Clk_period;
		Addr <=  "0010110010111";
		Trees_din <= x"0e003210";
		wait for Clk_period;
		Addr <=  "0010110011000";
		Trees_din <= x"16006d08";
		wait for Clk_period;
		Addr <=  "0010110011001";
		Trees_din <= x"16006004";
		wait for Clk_period;
		Addr <=  "0010110011010";
		Trees_din <= x"ffe0170d";
		wait for Clk_period;
		Addr <=  "0010110011011";
		Trees_din <= x"ff76170d";
		wait for Clk_period;
		Addr <=  "0010110011100";
		Trees_din <= x"16006d04";
		wait for Clk_period;
		Addr <=  "0010110011101";
		Trees_din <= x"0097170d";
		wait for Clk_period;
		Addr <=  "0010110011110";
		Trees_din <= x"ffdd170d";
		wait for Clk_period;
		Addr <=  "0010110011111";
		Trees_din <= x"16007408";
		wait for Clk_period;
		Addr <=  "0010110100000";
		Trees_din <= x"0009fa04";
		wait for Clk_period;
		Addr <=  "0010110100001";
		Trees_din <= x"007a170d";
		wait for Clk_period;
		Addr <=  "0010110100010";
		Trees_din <= x"ff9a170d";
		wait for Clk_period;
		Addr <=  "0010110100011";
		Trees_din <= x"1c028704";
		wait for Clk_period;
		Addr <=  "0010110100100";
		Trees_din <= x"ff99170d";
		wait for Clk_period;
		Addr <=  "0010110100101";
		Trees_din <= x"006a170d";
		wait for Clk_period;
		Addr <=  "0010110100110";
		Trees_din <= x"020b032c";
		wait for Clk_period;
		Addr <=  "0010110100111";
		Trees_din <= x"10004814";
		wait for Clk_period;
		Addr <=  "0010110101000";
		Trees_din <= x"0d008508";
		wait for Clk_period;
		Addr <=  "0010110101001";
		Trees_din <= x"1e025004";
		wait for Clk_period;
		Addr <=  "0010110101010";
		Trees_din <= x"0030170d";
		wait for Clk_period;
		Addr <=  "0010110101011";
		Trees_din <= x"ff84170d";
		wait for Clk_period;
		Addr <=  "0010110101100";
		Trees_din <= x"08004308";
		wait for Clk_period;
		Addr <=  "0010110101101";
		Trees_din <= x"03f82104";
		wait for Clk_period;
		Addr <=  "0010110101110";
		Trees_din <= x"0006170d";
		wait for Clk_period;
		Addr <=  "0010110101111";
		Trees_din <= x"0089170d";
		wait for Clk_period;
		Addr <=  "0010110110000";
		Trees_din <= x"ffd8170d";
		wait for Clk_period;
		Addr <=  "0010110110001";
		Trees_din <= x"000e8010";
		wait for Clk_period;
		Addr <=  "0010110110010";
		Trees_din <= x"05f4e008";
		wait for Clk_period;
		Addr <=  "0010110110011";
		Trees_din <= x"17f81704";
		wait for Clk_period;
		Addr <=  "0010110110100";
		Trees_din <= x"ffdf170d";
		wait for Clk_period;
		Addr <=  "0010110110101";
		Trees_din <= x"001f170d";
		wait for Clk_period;
		Addr <=  "0010110110110";
		Trees_din <= x"15004104";
		wait for Clk_period;
		Addr <=  "0010110110111";
		Trees_din <= x"001a170d";
		wait for Clk_period;
		Addr <=  "0010110111000";
		Trees_din <= x"008a170d";
		wait for Clk_period;
		Addr <=  "0010110111001";
		Trees_din <= x"08004204";
		wait for Clk_period;
		Addr <=  "0010110111010";
		Trees_din <= x"0040170d";
		wait for Clk_period;
		Addr <=  "0010110111011";
		Trees_din <= x"ffaa170d";
		wait for Clk_period;
		Addr <=  "0010110111100";
		Trees_din <= x"04057d04";
		wait for Clk_period;
		Addr <=  "0010110111101";
		Trees_din <= x"ff90170d";
		wait for Clk_period;
		Addr <=  "0010110111110";
		Trees_din <= x"1800d808";
		wait for Clk_period;
		Addr <=  "0010110111111";
		Trees_din <= x"03f7c704";
		wait for Clk_period;
		Addr <=  "0010111000000";
		Trees_din <= x"0006170d";
		wait for Clk_period;
		Addr <=  "0010111000001";
		Trees_din <= x"0066170d";
		wait for Clk_period;
		Addr <=  "0010111000010";
		Trees_din <= x"ffa4170d";
		wait for Clk_period;
		Addr <=  "0010111000011";
		Trees_din <= x"010e324c";
		wait for Clk_period;
		Addr <=  "0010111000100";
		Trees_din <= x"0400631c";
		wait for Clk_period;
		Addr <=  "0010111000101";
		Trees_din <= x"1403db08";
		wait for Clk_period;
		Addr <=  "0010111000110";
		Trees_din <= x"0a003d04";
		wait for Clk_period;
		Addr <=  "0010111000111";
		Trees_din <= x"fff117b9";
		wait for Clk_period;
		Addr <=  "0010111001000";
		Trees_din <= x"ff7e17b9";
		wait for Clk_period;
		Addr <=  "0010111001001";
		Trees_din <= x"02054608";
		wait for Clk_period;
		Addr <=  "0010111001010";
		Trees_din <= x"08003204";
		wait for Clk_period;
		Addr <=  "0010111001011";
		Trees_din <= x"000f17b9";
		wait for Clk_period;
		Addr <=  "0010111001100";
		Trees_din <= x"ff8817b9";
		wait for Clk_period;
		Addr <=  "0010111001101";
		Trees_din <= x"02074f08";
		wait for Clk_period;
		Addr <=  "0010111001110";
		Trees_din <= x"1403ff04";
		wait for Clk_period;
		Addr <=  "0010111001111";
		Trees_din <= x"00a217b9";
		wait for Clk_period;
		Addr <=  "0010111010000";
		Trees_din <= x"ffe517b9";
		wait for Clk_period;
		Addr <=  "0010111010001";
		Trees_din <= x"ff8e17b9";
		wait for Clk_period;
		Addr <=  "0010111010010";
		Trees_din <= x"06ff6f14";
		wait for Clk_period;
		Addr <=  "0010111010011";
		Trees_din <= x"10005510";
		wait for Clk_period;
		Addr <=  "0010111010100";
		Trees_din <= x"0207ba08";
		wait for Clk_period;
		Addr <=  "0010111010101";
		Trees_din <= x"03f9c504";
		wait for Clk_period;
		Addr <=  "0010111010110";
		Trees_din <= x"006c17b9";
		wait for Clk_period;
		Addr <=  "0010111010111";
		Trees_din <= x"ffd517b9";
		wait for Clk_period;
		Addr <=  "0010111011000";
		Trees_din <= x"0e003504";
		wait for Clk_period;
		Addr <=  "0010111011001";
		Trees_din <= x"ffa117b9";
		wait for Clk_period;
		Addr <=  "0010111011010";
		Trees_din <= x"002917b9";
		wait for Clk_period;
		Addr <=  "0010111011011";
		Trees_din <= x"ffa717b9";
		wait for Clk_period;
		Addr <=  "0010111011100";
		Trees_din <= x"04057d10";
		wait for Clk_period;
		Addr <=  "0010111011101";
		Trees_din <= x"0400b208";
		wait for Clk_period;
		Addr <=  "0010111011110";
		Trees_din <= x"05f55d04";
		wait for Clk_period;
		Addr <=  "0010111011111";
		Trees_din <= x"009f17b9";
		wait for Clk_period;
		Addr <=  "0010111100000";
		Trees_din <= x"000517b9";
		wait for Clk_period;
		Addr <=  "0010111100001";
		Trees_din <= x"010d5f04";
		wait for Clk_period;
		Addr <=  "0010111100010";
		Trees_din <= x"ffb517b9";
		wait for Clk_period;
		Addr <=  "0010111100011";
		Trees_din <= x"003917b9";
		wait for Clk_period;
		Addr <=  "0010111100100";
		Trees_din <= x"020d7908";
		wait for Clk_period;
		Addr <=  "0010111100101";
		Trees_din <= x"000f3604";
		wait for Clk_period;
		Addr <=  "0010111100110";
		Trees_din <= x"006017b9";
		wait for Clk_period;
		Addr <=  "0010111100111";
		Trees_din <= x"ffe117b9";
		wait for Clk_period;
		Addr <=  "0010111101000";
		Trees_din <= x"ffd017b9";
		wait for Clk_period;
		Addr <=  "0010111101001";
		Trees_din <= x"14016404";
		wait for Clk_period;
		Addr <=  "0010111101010";
		Trees_din <= x"003417b9";
		wait for Clk_period;
		Addr <=  "0010111101011";
		Trees_din <= x"05f22e04";
		wait for Clk_period;
		Addr <=  "0010111101100";
		Trees_din <= x"000817b9";
		wait for Clk_period;
		Addr <=  "0010111101101";
		Trees_din <= x"ff7a17b9";
		wait for Clk_period;
		Addr <=  "0010111101110";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  6
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"050b6020";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"0504f810";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"05009804";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"ff51004d";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"03fab204";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"ff5c004d";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"02029204";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"00df004d";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"ff8c004d";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"04fc450c";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"0107ec08";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"02021704";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"01b0004d";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"0037004d";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"ffa4004d";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"ff6d004d";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"02093404";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"047f004d";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"00ca004d";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"050b6020";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"0504f810";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"05009804";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"ff560099";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"03fab204";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"ff620099";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"1403fc04";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"ff8f0099";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"00bc0099";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"02003c08";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"1afc8e04";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"ffa20099";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"01bb0099";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"1b028404";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"ff700099";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"003c0099";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"1ef8ef04";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"00850099";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"01b00099";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"050b6020";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"0504f814";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"05009804";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"ff5a00fd";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"03fab204";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"ff6700fd";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"08003d08";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"0a004004";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"00d400fd";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"003000fd";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"ff8c00fd";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"1b028608";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"02fed204";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"007700fd";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"ff7200fd";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"00fa00fd";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"020b2110";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"2003fe04";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"004800fd";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"1a02ba08";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"00086304";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"013d00fd";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"006900fd";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"005c00fd";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"002500fd";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"050b6020";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"0504f814";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"05009804";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"ff5c0171";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"03fab204";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"ff6b0171";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"04fb1404";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"ff8f0171";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"05016304";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"00c70171";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"00220171";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"1e028608";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"02fed204";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"00630171";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"ff760171";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"00d40171";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"0a003a08";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"1b027a04";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"ffc90171";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"00ba0171";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"0511b810";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"1404000c";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"1e025204";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"fff00171";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"0900e604";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"010a0171";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"00540171";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"ffc20171";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"010b0171";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"050b6020";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"05009804";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"ff5e01dd";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"03fab20c";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"04f8d408";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"08004004";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"ff9f01dd";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"00ad01dd";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"ff6901dd";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"1b025604";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"ff9a01dd";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"15003404";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"ffa701dd";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"0c00a904";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"001201dd";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"012401dd";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"0511b810";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"0400030c";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"1e025204";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"ffe901dd";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"11002104";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"001301dd";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"00e201dd";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"ff7301dd";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"2003fe04";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"001c01dd";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"00e801dd";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"05075f14";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"05009804";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"ff600241";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"03fab204";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"ff6f0241";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"0105ce08";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"1101f804";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"ff7f0241";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"00830241";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"00cf0241";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"0511b818";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"04000314";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"08003908";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"03f9bb04";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"ff810241";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"00330241";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"0b006104";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"ffc40241";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"04f80e04";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"00070241";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"00cf0241";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"ff7a0241";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"2003fe04";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"00110241";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"00d20241";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"0504f810";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"05009804";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"ff6102b5";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"08003d08";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"08003a04";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"ff9302b5";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"00a602b5";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"ff7402b5";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"050b6010";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"14037208";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"0c00c404";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"00b902b5";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"ffef02b5";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"14040004";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"ff8602b5";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"001a02b5";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"0a003a08";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"12007804";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"ffa802b5";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"007b02b5";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"0511b810";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"0d000608";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"03f9bb04";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"ff6f02b5";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"006c02b5";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"17f73504";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"ffcb02b5";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"00b302b5";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"00c302b5";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"0504f810";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"05009804";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"ff620311";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"08003d08";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"08003a04";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"ff980311";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"008c0311";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"ff780311";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"0511b818";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"04000314";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"06039b0c";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"1e023304";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"ffe00311";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"0900d604";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"00b20311";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"00390311";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"0f004404";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"ff6c0311";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"00790311";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"ff7e0311";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"2003fe04";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"fff40311";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"00b90311";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"0504f810";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"05009804";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"ff630371";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"08003d08";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"08003a04";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"ff9e0371";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"00780371";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"ff7d0371";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"0511b818";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"04000314";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"0107ec10";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"06039b08";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"07fcb204";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"fff00371";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"009c0371";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"1e027d04";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"ff780371";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"00720371";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"ff9b0371";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"ff880371";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"2003fe04";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"ffec0371";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"00b10371";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"050b6018";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"05009804";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"ff6403d5";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"03fab208";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"1afd5404";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"ff7603d5";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"002003d5";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"0105ce08";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"1b027204";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"ff8903d5";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"006403d5";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"008403d5";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"0a003a08";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"1b027a04";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"ff9b03d5";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"005903d5";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"0511b810";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"08003c08";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"0a004504";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"006203d5";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"ff9603d5";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"06039b04";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"00a803d5";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"000b03d5";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"00ac03d5";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"0504f810";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"05009804";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"ff650441";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"0900e908";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"06fcca04";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"fff20441";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"ff830441";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"00340441";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"05145524";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"08003c10";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"03fb860c";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"0d000a04";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"ff660441";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"0d007004";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"00380441";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"ffb10441";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"00520441";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"1403e508";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"18032904";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"00a60441";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"00050441";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"08004104";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"00650441";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"07018c04";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"00130441";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"ff8c0441";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"00a70441";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"0504f810";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"05009804";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"ff650495";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"0a003e04";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"00320495";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"0d000904";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"fffb0495";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"ff860495";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"05145518";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"0a003e08";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"1101b804";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"ff850495";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"00020495";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"04008e0c";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"0d000604";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"ffe30495";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"050b6004";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"00210495";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"00980495";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"ff9d0495";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"00a20495";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"0504f810";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"05009804";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"ff6604f9";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"08003d08";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"08003a04";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"ffaf04f9";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"006204f9";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"ff8c04f9";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"05145520";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"1e027a14";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"06025d0c";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"1d027608";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"06fefa04";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"ffef04f9";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"007804f9";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"ff9704f9";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"04fc9604";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"ffd904f9";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"ff7504f9";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"0b008508";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"0f008104";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"002a04f9";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"009504f9";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"001204f9";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"009e04f9";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"0504f810";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"05009804";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"ff670565";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"03fab204";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"ff910565";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"0d006104";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"ffdd0565";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"004e0565";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"05145524";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"08003c10";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"03fb860c";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"0d000a04";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"ff760565";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"17f82904";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"000f0565";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"ffd40565";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"003d0565";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"1403e508";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"11028f04";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"00890565";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"000e0565";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"08004104";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"00520565";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"0900b804";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"00070565";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"ff9b0565";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"009a0565";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"050b6014";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"05009804";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"ff6705b1";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"01056008";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"03fee004";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"ff7f05b1";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"000d05b1";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"1afc9604";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"ffdb05b1";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"007005b1";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"0a003a04";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"ffd205b1";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"0511b80c";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"1e025204";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"ffc105b1";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"08003a04";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"ffed05b1";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"007d05b1";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"009805b1";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"050b6014";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"05009804";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"ff6805fd";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"01056008";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"03fee004";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"ff8305fd";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"000a05fd";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"1afc9604";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"ffde05fd";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"006805fd";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"0a003a04";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"ffd205fd";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"0511b80c";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"0c00b308";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"0b007304";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"003c05fd";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"ff9f05fd";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"007c05fd";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"009405fd";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"05075f14";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"05009804";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"ff68065d";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"03fab204";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"ff95065d";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"03fbd204";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"005d065d";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"1b026b04";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"ff9d065d";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"002c065d";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"05145518";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"1e027a10";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"06025d0c";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"1d027508";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"0a004504";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"006a065d";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"ffff065d";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"ffaa065d";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"ff94065d";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"0e002904";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"001d065d";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"007b065d";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"008f065d";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"050b6014";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"05009804";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"ff6906a1";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"01056008";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"03fee004";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"ff8906a1";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"000406a1";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"1afc9804";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"ffe006a1";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"005806a1";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"0a003a04";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"ffce06a1";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"1e025204";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"000206a1";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"14040004";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"008a06a1";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"000806a1";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"05009804";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"ff6a06e5";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"0514551c";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"0d002208";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"06ffe304";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"001206e5";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"ff9106e5";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"050b600c";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"1b026804";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"ffaf06e5";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"03fab204";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"ffdb06e5";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"005106e5";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"0c00a404";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"000006e5";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"007606e5";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"008706e5";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"05009804";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"ff6b0731";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"05145520";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"1e027b14";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"06025d10";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"18005208";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"02037e04";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"00610731";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"ffe40731";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"0c00af04";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"ff9a0731";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"00230731";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"ff910731";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"05075f04";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"ffdc0731";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"19000104";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"001d0731";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"006c0731";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"00830731";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"05009804";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"ff6c0775";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"0514551c";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"0d002208";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"06ffe304";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"000b0775";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"ffa00775";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"050b600c";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"1b026804";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"ffb80775";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"03fab204";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"ffe00775";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"004b0775";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"0c00a404";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"00050775";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"006c0775";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"007f0775";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"05009804";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"ff6d07b9";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"0514551c";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"08003a08";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"00006604";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"fffd07b9";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"ffa207b9";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"0c00a808";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"00ffa604";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"002f07b9";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"ffac07b9";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"06fe8904";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"fff407b9";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"1afc1004";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"001507b9";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"006407b9";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"007b07b9";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"05009804";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"ff6e07fd";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"0514551c";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"0d002208";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"03f9bb04";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"ffa907fd";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"000a07fd";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"050b600c";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"02003c04";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"002d07fd";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"0d007404";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"001807fd";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"ff9c07fd";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"0c00a404";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"000f07fd";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"006507fd";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"007807fd";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"0504f80c";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"05009804";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"ff6f0841";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"08003d04";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"00180841";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"ffab0841";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"05145514";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"0a003e04";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"ffb90841";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"0e002e08";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"0c00b304";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"ffb40841";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"00310841";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"17f7d704";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"00150841";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"005f0841";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"00740841";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"05075f10";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"05009804";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"ff710885";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"0105e908";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"0b006904";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"fff90885";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"ffa30885";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"00190885";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"0a003e04";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"ffdf0885";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"0511b80c";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"08003d04";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"ffd70885";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"04fc7e04";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"005a0885";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"00100885";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"00730885";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"05009804";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"ff7308c1";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"05145518";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"0d002208";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"06ffe304";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"000708c1";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"ffb108c1";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"050b6008";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"03fab204";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"ffc008c1";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"001608c1";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"0c00a404";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"000e08c1";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"005c08c1";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"006c08c1";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  7
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"02089668";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"02069e2c";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"010eef20";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"0203d810";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"2003ff08";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"03f94e04";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"ff840185";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"00ca0185";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"04f77004";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"ffcb0185";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"ff610185";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"000ba108";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"08004304";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"ffb60185";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"000f0185";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"0e005304";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"ff5e0185";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"00370185";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"22002004";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"ff570185";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"00093304";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"ff900185";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"00370185";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"07fdaf20";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"000cc010";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"010e5008";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"04000304";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"ffd70185";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"00a50185";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"04003a04";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"ff570185";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"ffa10185";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"0405f108";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"06fbe104";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"ffe80185";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"ff590185";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"00110d04";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"005b0185";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"ff700185";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"0300dc10";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"000b1d08";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"02079004";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"00a30185";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"022d0185";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"08003104";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"00370185";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"ff680185";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"0a005008";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"05fa8504";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"ff5d0185";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"00370185";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"012b0185";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"000cc030";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"03122d20";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"010bfd10";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"060d0408";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"020b0304";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"02250185";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"03a80185";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"02107804";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"000e0185";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"022f0185";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"06fe5208";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"12007804";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"022f0185";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"ffa40185";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"02091004";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"009f0185";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"ff830185";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"17fff90c";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"07fd7a08";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"01004904";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"00370185";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"ff9c0185";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"ff5b0185";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"00370185";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"0010c51c";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"020b2110";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"07f62508";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"0c00a904";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"01b00185";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"ff9c0185";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"11014804";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"ff620185";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"00260185";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"03f74208";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"12008604";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"02bc0185";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"00210185";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"ff8c0185";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"1e02870c";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"03f8e608";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"13040004";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"ff550185";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"00000185";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"000f0185";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"00890185";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"02081960";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"010e503c";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"02061a1c";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"0203420c";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"1cfd6504";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"004002f1";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"19000a04";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"ff5e02f1";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"ffa702f1";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"000ba108";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"21000004";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"ffc602f1";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"005202f1";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"12009d04";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"ff5902f1";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"000702f1";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"000be510";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"16003e08";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"0007b504";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"022b02f1";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"002d02f1";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"030c2c04";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"004402f1";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"ff6402f1";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"0c00a408";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"0c009f04";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"ff7002f1";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"008d02f1";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"03fa5204";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"ff5b02f1";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"000302f1";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"0207c518";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"22002010";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"0a005c08";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"0a004304";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"ff6e02f1";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"ff5702f1";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"05f45704";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"ff8d02f1";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"004002f1";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"0c00bb04";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"ff9902f1";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"003a02f1";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"0b007a04";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"ff7502f1";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"06ff5b04";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"ffa902f1";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"00db02f1";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"000e8030";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"03122d20";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"010cb710";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"04098208";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"020a8004";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"00fb02f1";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"018b02f1";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"16005f04";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"002b02f1";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"ff5c02f1";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"15004108";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"06fc4b04";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"00c702f1";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"ff7602f1";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"0f000404";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"ff8002f1";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"01b302f1";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"1b04820c";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"020b5c04";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"ff6102f1";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"0b006d04";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"003e02f1";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"ff9002f1";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"003502f1";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"0010c518";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"0405aa10";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"15004708";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"16005d04";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"001402f1";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"ff6602f1";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"08004504";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"ff9b02f1";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"011d02f1";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"1101b804";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"019d02f1";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"000d02f1";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"1f02870c";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"0a003e08";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"17f78404";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"00b302f1";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"ff7802f1";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"ff5b02f1";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"005a02f1";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"0208195c";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"010e5040";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"02069620";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"0203d810";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"11000008";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"0202f304";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"ff9a043d";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"00cf043d";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"0d027304";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"ff6c043d";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"ffd1043d";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"000ba108";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"12008704";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"ffd4043d";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"0057043d";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"15005204";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"ff68043d";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"0039043d";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"000cc010";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"00003a08";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"0a004e04";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"ff66043d";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"00af043d";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"14034d04";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"ffd0043d";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"007b043d";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"06fd4908";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"05f42904";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"0094043d";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"ff83043d";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"0a003b04";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"0020043d";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"ff5f043d";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"0207c514";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"2200200c";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"05f4c304";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"ff5f043d";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"000b3304";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"ff6d043d";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"fff0043d";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"0b008404";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"0044043d";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"ffa0043d";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"1800e104";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"ff7b043d";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"005f043d";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"000fa830";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"03122d20";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"010cb710";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"000ac708";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"06112304";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"0101043d";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"ffc0043d";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"020eae04";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"0055043d";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"0169043d";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"15004208";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"06fc4b04";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"00b3043d";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"ff7b043d";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"0f000404";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"ff83043d";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"0141043d";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"1b04820c";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"00fc1108";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"0d00c504";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"0042043d";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"ff9e043d";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"ff66043d";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"0032043d";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"1b024908";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"03f60504";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"ff88043d";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"012c043d";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"07fbf108";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"07f39d04";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"fff6043d";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"ff5e043d";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"12007704";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"ff81043d";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"0c00c304";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"0119043d";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"ffa8043d";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"0207ad64";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"010e5038";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"0203d818";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"2003ff08";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"03f87604";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"ff9d0599";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"00d30599";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"0b005a08";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"0e004404";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"00d50599";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"ff870599";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"04f77004";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"00030599";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"ff720599";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"000be510";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"01ff1108";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"0b008a04";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"ff620599";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"00310599";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"010c1204";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"00300599";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"ffcf0599";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"03fa5208";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"0203f204";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"00400599";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"ff770599";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"07f7e704";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"00c40599";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"ff8a0599";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"0a004320";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"20040010";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"06fcca08";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"07ffc304";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"010a0599";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"ff920599";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"02061004";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"ff6d0599";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"00290599";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"010e8408";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"07f93504";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"00470599";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"ff960599";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"0b008e04";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"ff6c0599";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"ffcc0599";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"0a005c04";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"ff5e0599";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"0e002604";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"ff9e0599";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"00420599";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"000fa82c";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"03145b20";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"020a8010";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"04032308";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"06099f04";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"008e0599";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"ff7b0599";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"1801fb04";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"ff5b0599";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"00420599";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"040a8408";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"14022704";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"000a0599";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"00d70599";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"0900c504";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"ff600599";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"008f0599";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"0900eb04";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"ff690599";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"15003d04";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"00420599";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"ffa80599";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"05f53b08";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"11000804";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"00240599";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"ff630599";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"15003910";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"0c00b808";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"0900e304";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"01960599";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"00360599";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"03f1e204";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"003a0599";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"ff870599";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"0b008104";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"ff6d0599";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"003d0599";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"02076e4c";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"010eef34";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"02034214";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"0d02790c";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"08001d04";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"004306ed";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"04f68e04";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"003a06ed";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"ff6a06ed";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"04f9f604";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"00ee06ed";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"ff7606ed";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"0006ee10";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"00042c08";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"0a003c04";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"00db06ed";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"ffcd06ed";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"06ff3f04";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"00b806ed";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"001006ed";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"03fc1e08";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"07fcca04";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"ff8e06ed";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"ffd006ed";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"0008d204";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"ff8206ed";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"018506ed";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"22002014";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"05f4c304";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"ff6406ed";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"0205c008";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"000b3304";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"ff6c06ed";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"ffe406ed";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"03f84004";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"00d706ed";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"ff8006ed";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"000c06ed";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"000ce328";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"03145b20";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"010bdd10";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"0d003908";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"0e005304";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"00bd06ed";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"ff7106ed";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"020e3704";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"004c06ed";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"00da06ed";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"0d007d08";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"0b006204";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"011206ed";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"ff8306ed";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"0a004204";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"ffc406ed";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"00d406ed";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"00fc1104";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"fffc06ed";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"ff6d06ed";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"020a0018";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"06fc0308";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"0900df04";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"ffa806ed";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"00d206ed";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"19000408";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"05f74304";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"ff6106ed";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"001c06ed";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"19000504";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"00d206ed";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"ffa306ed";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"01079710";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"020e3708";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"0a004f04";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"ff6d06ed";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"005d06ed";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"0010c504";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"00de06ed";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"ff9e06ed";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"03f4a508";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"1100a204";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"00b706ed";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"ffa206ed";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"08003304";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"002b06ed";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"018006ed";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"02076e48";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"010eef30";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"0203d814";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"2003fe04";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"005307e9";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"0b005a08";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"0f000604";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"ff9107e9";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"00dc07e9";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"04f77004";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"001407e9";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"ff7c07e9";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"000ba110";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"12009f08";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"01ff1104";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"ff6707e9";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"000707e9";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"1801b004";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"01c907e9";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"ffa207e9";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"08004004";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"ff6507e9";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"08004104";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"009107e9";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"ffa207e9";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"22002014";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"05f4c304";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"ff6707e9";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"0205c008";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"000b3304";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"ff7107e9";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"ffee07e9";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"0900e104";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"ff8607e9";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"00c307e9";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"001507e9";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"0011792c";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"020f5a1c";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"00fe5f10";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"0b009408";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"00fc1104";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"fffc07e9";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"ff5c07e9";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"01036904";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"000e07e9";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"00a607e9";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"010ff908";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"04032304";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"006807e9";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"000107e9";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"ff6d07e9";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"00fe1808";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"0f002704";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"ffbb07e9";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"00a007e9";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"14040004";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"00e507e9";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"002907e9";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"1f028708";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"17f71304";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"001b07e9";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"ff6807e9";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"007307e9";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"0206dd58";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"010c8438";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"02034218";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"0d027910";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"19001b08";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"03f60e04";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"ffb40955";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"ff650955";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"0108b504";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"ff8f0955";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"00c20955";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"04f9f604";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"01250955";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"ff890955";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"000b1d10";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"0e003808";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"08004404";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"00090955";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"00fb0955";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"11000604";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"00860955";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"ffb40955";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"05f2e408";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"0f000704";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"00db0955";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"ff9d0955";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"12008904";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"ff660955";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"00150955";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"0a004614";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"01119e10";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"16007c08";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"12008904";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"ff9b0955";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"00540955";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"05f59f04";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"ffbe0955";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"012e0955";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"ff680955";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"0a005c04";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"ff620955";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"1f026704";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"ffa70955";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"00470955";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"0209bd3c";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"04022520";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"0605ab10";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"17fdec08";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"03fb1b04";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"00590955";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"fff30955";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"1e061a04";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"ff550955";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"00370955";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"08003708";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"07fd3804";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"ff9d0955";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"01270955";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"04fb7f04";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"005b0955";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"ff4c0955";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"03f98410";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"0405f108";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"0a003d04";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"00280955";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"ff560955";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"0f001004";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"ff7b0955";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"005f0955";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"09009704";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"01390955";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"0d00d604";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"ff7f0955";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"003e0955";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"0015b320";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"00ff6310";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"0608d708";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"020b2104";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"ffa00955";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"00830955";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"01f76404";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"00170955";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"ff520955";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"040a8408";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"0d005f04";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"00960955";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"00530955";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"0900c804";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"ff650955";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"004d0955";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"ff7c0955";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"02088c54";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"010eef38";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"000bff20";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"02034210";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"19000a08";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"0008a904";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"ff6f0a85";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"00160a85";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"0f003204";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"010e0a85";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"ffa10a85";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"12008608";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"16008104";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"ffe40a85";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"00490a85";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"03f95504";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"fff70a85";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"00a90a85";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"02061a08";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"0c00ef04";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"ff670a85";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"00310a85";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"0900c108";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"06fd8f04";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"003f0a85";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"ff650a85";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"0d01de04";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"ffca0a85";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"00e50a85";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"0a004314";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"0a004310";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"20040008";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"05f51e04";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"ffaf0a85";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"00aa0a85";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"14040004";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"ff7c0a85";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"00150a85";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"00850a85";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"13009f04";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"00360a85";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"ff660a85";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"0210783c";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"0104dc20";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"0008c210";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"10004408";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"16006304";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"00220a85";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"ff4c0a85";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"10004c04";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"00a90a85";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"00190a85";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"1f026908";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"0d00da04";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"ff500a85";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"002b0a85";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"1b026a04";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"00d90a85";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"fffc0a85";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"15004e10";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"0c00ae08";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"14036004";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"00090a85";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"00a50a85";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"07f97504";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"ffbb0a85";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"00740a85";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"07ff4308";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"16009604";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"00130a85";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"ff430a85";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"00bc0a85";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"06112304";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"00c40a85";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"ffef0a85";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"02058658";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"010c1230";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"010b131c";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"21000610";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"0c007008";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"15004a04";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"00c00bf9";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"ff9e0bf9";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"11032604";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"ff9d0bf9";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"00860bf9";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"05f70f04";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"ff910bf9";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"22000104";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"00cf0bf9";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"ffa90bf9";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"0c00a608";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"06fd3704";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"00430bf9";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"ff890bf9";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"0203d104";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"ffa00bf9";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"1403e804";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"00350bf9";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"02800bf9";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"0c00e81c";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"0900e90c";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"10003404";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"002f0bf9";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"19002c04";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"ff6e0bf9";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"ffe00bf9";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"0900eb08";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"04fd5404";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"ffa50bf9";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"01760bf9";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"0a003d04";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"00490bf9";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"ff700bf9";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"010d0204";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"01110bf9";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"08003f04";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"ff860bf9";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"00440bf9";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"0209ee3c";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"04022520";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"000cc010";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"0605ab08";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"03103e04";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"00390bf9";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"ff720bf9";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"08003704";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"00630bf9";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"ff7e0bf9";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"04017708";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"0f000104";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"004b0bf9";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"ff650bf9";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"1403ef04";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"01410bf9";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"ff910bf9";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"03f98410";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"0d017008";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"01f6a404";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"00130bf9";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"ff660bf9";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"0d020504";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"007a0bf9";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"ff7c0bf9";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"1b025c04";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"ff790bf9";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"0404a704";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"00dd0bf9";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"ff9c0bf9";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"02107820";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"0103ef10";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"05f57d08";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"07024804";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"ff7b0bf9";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"00970bf9";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"10004404";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"ffeb0bf9";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"00530bf9";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"0d00ad08";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"15002904";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"ff4d0bf9";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"008c0bf9";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"1c028704";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"00100bf9";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"01110bf9";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"06112304";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"00b60bf9";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"fff00bf9";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"02058640";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"12008724";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"000b4520";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"04fc6810";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"00fc6608";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"0a003f04";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"00bb0cdd";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"ff9e0cdd";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"13040004";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"ff7a0cdd";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"002a0cdd";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"0900e408";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"19002104";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"ffaf0cdd";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"00b20cdd";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"0008a904";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"ffe00cdd";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"01120cdd";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"ff680cdd";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"0a004d18";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"0e001f08";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"003b0cdd";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"ff7b0cdd";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"0b008308";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"04ff7404";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"ff900cdd";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"00310cdd";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"02048604";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"017f0cdd";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"ffef0cdd";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"ff6e0cdd";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"020f5a24";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"010ff918";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"00120e10";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"10004408";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"010a1304";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"00220cdd";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"ffcf0cdd";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"1302e104";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"fffd0cdd";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"00480cdd";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"1f028704";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"ff700cdd";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"006e0cdd";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"05f55d08";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"0b006004";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"00210cdd";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"ff6d0cdd";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"00490cdd";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"00fe1808";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"0f002704";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"ffbf0cdd";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"00640cdd";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"14040004";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"00ac0cdd";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"fff50cdd";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"02058654";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"010c1230";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"010b131c";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"0800440c";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"10004204";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"ff650e21";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"1afc8504";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"00340e21";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"ff850e21";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"0e003608";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"19001104";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"01040e21";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"ff8f0e21";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"13040004";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"ff690e21";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"00f10e21";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"0c00a608";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"13037804";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"00440e21";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"ff960e21";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"0203d104";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"ffa90e21";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"08003e04";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"005a0e21";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"019a0e21";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"0c00e818";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"0900e90c";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"15002c04";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"003e0e21";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"02056b04";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"ff750e21";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"00010e21";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"06fd9a08";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"04fcc104";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"ff8c0e21";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"01020e21";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"ff780e21";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"0e002308";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"00390e21";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"ff920e21";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"00c00e21";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"020f5a40";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"04fdd620";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"03f61810";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"1403fc08";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"0f002c04";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"018b0e21";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"00420e21";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"12007304";
		wait for Clk_period;
		Addr <=  "0001101101001";
		Trees_din <= x"00490e21";
		wait for Clk_period;
		Addr <=  "0001101101010";
		Trees_din <= x"ff830e21";
		wait for Clk_period;
		Addr <=  "0001101101011";
		Trees_din <= x"0f010808";
		wait for Clk_period;
		Addr <=  "0001101101100";
		Trees_din <= x"0a004504";
		wait for Clk_period;
		Addr <=  "0001101101101";
		Trees_din <= x"ffdf0e21";
		wait for Clk_period;
		Addr <=  "0001101101110";
		Trees_din <= x"004e0e21";
		wait for Clk_period;
		Addr <=  "0001101101111";
		Trees_din <= x"010b3c04";
		wait for Clk_period;
		Addr <=  "0001101110000";
		Trees_din <= x"00c30e21";
		wait for Clk_period;
		Addr <=  "0001101110001";
		Trees_din <= x"ff820e21";
		wait for Clk_period;
		Addr <=  "0001101110010";
		Trees_din <= x"06fde610";
		wait for Clk_period;
		Addr <=  "0001101110011";
		Trees_din <= x"0c00ae08";
		wait for Clk_period;
		Addr <=  "0001101110100";
		Trees_din <= x"0c009604";
		wait for Clk_period;
		Addr <=  "0001101110101";
		Trees_din <= x"00060e21";
		wait for Clk_period;
		Addr <=  "0001101110110";
		Trees_din <= x"00fb0e21";
		wait for Clk_period;
		Addr <=  "0001101110111";
		Trees_din <= x"020a0004";
		wait for Clk_period;
		Addr <=  "0001101111000";
		Trees_din <= x"ff990e21";
		wait for Clk_period;
		Addr <=  "0001101111001";
		Trees_din <= x"008e0e21";
		wait for Clk_period;
		Addr <=  "0001101111010";
		Trees_din <= x"14035308";
		wait for Clk_period;
		Addr <=  "0001101111011";
		Trees_din <= x"02093404";
		wait for Clk_period;
		Addr <=  "0001101111100";
		Trees_din <= x"ff800e21";
		wait for Clk_period;
		Addr <=  "0001101111101";
		Trees_din <= x"fffe0e21";
		wait for Clk_period;
		Addr <=  "0001101111110";
		Trees_din <= x"01044d04";
		wait for Clk_period;
		Addr <=  "0001101111111";
		Trees_din <= x"ffd20e21";
		wait for Clk_period;
		Addr <=  "0001110000000";
		Trees_din <= x"001d0e21";
		wait for Clk_period;
		Addr <=  "0001110000001";
		Trees_din <= x"1404000c";
		wait for Clk_period;
		Addr <=  "0001110000010";
		Trees_din <= x"00fe1808";
		wait for Clk_period;
		Addr <=  "0001110000011";
		Trees_din <= x"08004004";
		wait for Clk_period;
		Addr <=  "0001110000100";
		Trees_din <= x"00310e21";
		wait for Clk_period;
		Addr <=  "0001110000101";
		Trees_din <= x"ffe20e21";
		wait for Clk_period;
		Addr <=  "0001110000110";
		Trees_din <= x"00a10e21";
		wait for Clk_period;
		Addr <=  "0001110000111";
		Trees_din <= x"fff00e21";
		wait for Clk_period;
		Addr <=  "0001110001000";
		Trees_din <= x"02088c4c";
		wait for Clk_period;
		Addr <=  "0001110001001";
		Trees_din <= x"05f4c32c";
		wait for Clk_period;
		Addr <=  "0001110001010";
		Trees_din <= x"010c2418";
		wait for Clk_period;
		Addr <=  "0001110001011";
		Trees_din <= x"13030908";
		wait for Clk_period;
		Addr <=  "0001110001100";
		Trees_din <= x"17f79d04";
		wait for Clk_period;
		Addr <=  "0001110001101";
		Trees_din <= x"001e0f7d";
		wait for Clk_period;
		Addr <=  "0001110001110";
		Trees_din <= x"ff670f7d";
		wait for Clk_period;
		Addr <=  "0001110001111";
		Trees_din <= x"0a003f08";
		wait for Clk_period;
		Addr <=  "0001110010000";
		Trees_din <= x"12008804";
		wait for Clk_period;
		Addr <=  "0001110010001";
		Trees_din <= x"ff640f7d";
		wait for Clk_period;
		Addr <=  "0001110010010";
		Trees_din <= x"000a0f7d";
		wait for Clk_period;
		Addr <=  "0001110010011";
		Trees_din <= x"11006f04";
		wait for Clk_period;
		Addr <=  "0001110010100";
		Trees_din <= x"ffb40f7d";
		wait for Clk_period;
		Addr <=  "0001110010101";
		Trees_din <= x"00860f7d";
		wait for Clk_period;
		Addr <=  "0001110010110";
		Trees_din <= x"1300e904";
		wait for Clk_period;
		Addr <=  "0001110010111";
		Trees_din <= x"005a0f7d";
		wait for Clk_period;
		Addr <=  "0001110011000";
		Trees_din <= x"06fde608";
		wait for Clk_period;
		Addr <=  "0001110011001";
		Trees_din <= x"02075704";
		wait for Clk_period;
		Addr <=  "0001110011010";
		Trees_din <= x"ff9e0f7d";
		wait for Clk_period;
		Addr <=  "0001110011011";
		Trees_din <= x"00900f7d";
		wait for Clk_period;
		Addr <=  "0001110011100";
		Trees_din <= x"05f2f604";
		wait for Clk_period;
		Addr <=  "0001110011101";
		Trees_din <= x"ffa60f7d";
		wait for Clk_period;
		Addr <=  "0001110011110";
		Trees_din <= x"ff650f7d";
		wait for Clk_period;
		Addr <=  "0001110011111";
		Trees_din <= x"05f4cf0c";
		wait for Clk_period;
		Addr <=  "0001110100000";
		Trees_din <= x"08004008";
		wait for Clk_period;
		Addr <=  "0001110100001";
		Trees_din <= x"010ab104";
		wait for Clk_period;
		Addr <=  "0001110100010";
		Trees_din <= x"00a60f7d";
		wait for Clk_period;
		Addr <=  "0001110100011";
		Trees_din <= x"ffa60f7d";
		wait for Clk_period;
		Addr <=  "0001110100100";
		Trees_din <= x"01f40f7d";
		wait for Clk_period;
		Addr <=  "0001110100101";
		Trees_din <= x"0200ea04";
		wait for Clk_period;
		Addr <=  "0001110100110";
		Trees_din <= x"ff710f7d";
		wait for Clk_period;
		Addr <=  "0001110100111";
		Trees_din <= x"1d026108";
		wait for Clk_period;
		Addr <=  "0001110101000";
		Trees_din <= x"1b025504";
		wait for Clk_period;
		Addr <=  "0001110101001";
		Trees_din <= x"00060f7d";
		wait for Clk_period;
		Addr <=  "0001110101010";
		Trees_din <= x"ffaa0f7d";
		wait for Clk_period;
		Addr <=  "0001110101011";
		Trees_din <= x"0006b204";
		wait for Clk_period;
		Addr <=  "0001110101100";
		Trees_din <= x"003a0f7d";
		wait for Clk_period;
		Addr <=  "0001110101101";
		Trees_din <= x"ffed0f7d";
		wait for Clk_period;
		Addr <=  "0001110101110";
		Trees_din <= x"0d001838";
		wait for Clk_period;
		Addr <=  "0001110101111";
		Trees_din <= x"10004e18";
		wait for Clk_period;
		Addr <=  "0001110110000";
		Trees_din <= x"04067d10";
		wait for Clk_period;
		Addr <=  "0001110110001";
		Trees_din <= x"06099f08";
		wait for Clk_period;
		Addr <=  "0001110110010";
		Trees_din <= x"030e8404";
		wait for Clk_period;
		Addr <=  "0001110110011";
		Trees_din <= x"00aa0f7d";
		wait for Clk_period;
		Addr <=  "0001110110100";
		Trees_din <= x"ff9e0f7d";
		wait for Clk_period;
		Addr <=  "0001110110101";
		Trees_din <= x"10004804";
		wait for Clk_period;
		Addr <=  "0001110110110";
		Trees_din <= x"ff530f7d";
		wait for Clk_period;
		Addr <=  "0001110110111";
		Trees_din <= x"008e0f7d";
		wait for Clk_period;
		Addr <=  "0001110111000";
		Trees_din <= x"0f00bc04";
		wait for Clk_period;
		Addr <=  "0001110111001";
		Trees_din <= x"ff4b0f7d";
		wait for Clk_period;
		Addr <=  "0001110111010";
		Trees_din <= x"004f0f7d";
		wait for Clk_period;
		Addr <=  "0001110111011";
		Trees_din <= x"00079110";
		wait for Clk_period;
		Addr <=  "0001110111100";
		Trees_din <= x"03f78d08";
		wait for Clk_period;
		Addr <=  "0001110111101";
		Trees_din <= x"0400a804";
		wait for Clk_period;
		Addr <=  "0001110111110";
		Trees_din <= x"ff6a0f7d";
		wait for Clk_period;
		Addr <=  "0001110111111";
		Trees_din <= x"00680f7d";
		wait for Clk_period;
		Addr <=  "0001111000000";
		Trees_din <= x"0003e304";
		wait for Clk_period;
		Addr <=  "0001111000001";
		Trees_din <= x"00180f7d";
		wait for Clk_period;
		Addr <=  "0001111000010";
		Trees_din <= x"00b90f7d";
		wait for Clk_period;
		Addr <=  "0001111000011";
		Trees_din <= x"07f79c08";
		wait for Clk_period;
		Addr <=  "0001111000100";
		Trees_din <= x"17f74c04";
		wait for Clk_period;
		Addr <=  "0001111000101";
		Trees_din <= x"ffe30f7d";
		wait for Clk_period;
		Addr <=  "0001111000110";
		Trees_din <= x"00b70f7d";
		wait for Clk_period;
		Addr <=  "0001111000111";
		Trees_din <= x"0e002704";
		wait for Clk_period;
		Addr <=  "0001111001000";
		Trees_din <= x"008f0f7d";
		wait for Clk_period;
		Addr <=  "0001111001001";
		Trees_din <= x"ff3e0f7d";
		wait for Clk_period;
		Addr <=  "0001111001010";
		Trees_din <= x"020e3718";
		wait for Clk_period;
		Addr <=  "0001111001011";
		Trees_din <= x"08004d10";
		wait for Clk_period;
		Addr <=  "0001111001100";
		Trees_din <= x"10004508";
		wait for Clk_period;
		Addr <=  "0001111001101";
		Trees_din <= x"0e002604";
		wait for Clk_period;
		Addr <=  "0001111001110";
		Trees_din <= x"00360f7d";
		wait for Clk_period;
		Addr <=  "0001111001111";
		Trees_din <= x"ffbf0f7d";
		wait for Clk_period;
		Addr <=  "0001111010000";
		Trees_din <= x"1afcbe04";
		wait for Clk_period;
		Addr <=  "0001111010001";
		Trees_din <= x"004f0f7d";
		wait for Clk_period;
		Addr <=  "0001111010010";
		Trees_din <= x"fff70f7d";
		wait for Clk_period;
		Addr <=  "0001111010011";
		Trees_din <= x"07fecd04";
		wait for Clk_period;
		Addr <=  "0001111010100";
		Trees_din <= x"ff140f7d";
		wait for Clk_period;
		Addr <=  "0001111010101";
		Trees_din <= x"00500f7d";
		wait for Clk_period;
		Addr <=  "0001111010110";
		Trees_din <= x"0611230c";
		wait for Clk_period;
		Addr <=  "0001111010111";
		Trees_din <= x"0e002f04";
		wait for Clk_period;
		Addr <=  "0001111011000";
		Trees_din <= x"00be0f7d";
		wait for Clk_period;
		Addr <=  "0001111011001";
		Trees_din <= x"1b025304";
		wait for Clk_period;
		Addr <=  "0001111011010";
		Trees_din <= x"ff6d0f7d";
		wait for Clk_period;
		Addr <=  "0001111011011";
		Trees_din <= x"00780f7d";
		wait for Clk_period;
		Addr <=  "0001111011100";
		Trees_din <= x"05f7db04";
		wait for Clk_period;
		Addr <=  "0001111011101";
		Trees_din <= x"00190f7d";
		wait for Clk_period;
		Addr <=  "0001111011110";
		Trees_din <= x"ffa10f7d";
		wait for Clk_period;
		Addr <=  "0001111011111";
		Trees_din <= x"02058648";
		wait for Clk_period;
		Addr <=  "0001111100000";
		Trees_din <= x"03f5f508";
		wait for Clk_period;
		Addr <=  "0001111100001";
		Trees_din <= x"00feb504";
		wait for Clk_period;
		Addr <=  "0001111100010";
		Trees_din <= x"00331091";
		wait for Clk_period;
		Addr <=  "0001111100011";
		Trees_din <= x"ff6b1091";
		wait for Clk_period;
		Addr <=  "0001111100100";
		Trees_din <= x"16006620";
		wait for Clk_period;
		Addr <=  "0001111100101";
		Trees_din <= x"08003e10";
		wait for Clk_period;
		Addr <=  "0001111100110";
		Trees_din <= x"18020208";
		wait for Clk_period;
		Addr <=  "0001111100111";
		Trees_din <= x"06014f04";
		wait for Clk_period;
		Addr <=  "0001111101000";
		Trees_din <= x"ff951091";
		wait for Clk_period;
		Addr <=  "0001111101001";
		Trees_din <= x"00271091";
		wait for Clk_period;
		Addr <=  "0001111101010";
		Trees_din <= x"19000104";
		wait for Clk_period;
		Addr <=  "0001111101011";
		Trees_din <= x"01131091";
		wait for Clk_period;
		Addr <=  "0001111101100";
		Trees_din <= x"ffa91091";
		wait for Clk_period;
		Addr <=  "0001111101101";
		Trees_din <= x"1403fe08";
		wait for Clk_period;
		Addr <=  "0001111101110";
		Trees_din <= x"1302c404";
		wait for Clk_period;
		Addr <=  "0001111101111";
		Trees_din <= x"00ba1091";
		wait for Clk_period;
		Addr <=  "0001111110000";
		Trees_din <= x"ffe71091";
		wait for Clk_period;
		Addr <=  "0001111110001";
		Trees_din <= x"04fe1e04";
		wait for Clk_period;
		Addr <=  "0001111110010";
		Trees_din <= x"00051091";
		wait for Clk_period;
		Addr <=  "0001111110011";
		Trees_din <= x"01bd1091";
		wait for Clk_period;
		Addr <=  "0001111110100";
		Trees_din <= x"0b006510";
		wait for Clk_period;
		Addr <=  "0001111110101";
		Trees_din <= x"08004108";
		wait for Clk_period;
		Addr <=  "0001111110110";
		Trees_din <= x"1afcf104";
		wait for Clk_period;
		Addr <=  "0001111110111";
		Trees_din <= x"016e1091";
		wait for Clk_period;
		Addr <=  "0001111111000";
		Trees_din <= x"ff861091";
		wait for Clk_period;
		Addr <=  "0001111111001";
		Trees_din <= x"01008904";
		wait for Clk_period;
		Addr <=  "0001111111010";
		Trees_din <= x"00281091";
		wait for Clk_period;
		Addr <=  "0001111111011";
		Trees_din <= x"ff731091";
		wait for Clk_period;
		Addr <=  "0001111111100";
		Trees_din <= x"0c007208";
		wait for Clk_period;
		Addr <=  "0001111111101";
		Trees_din <= x"04fc7604";
		wait for Clk_period;
		Addr <=  "0001111111110";
		Trees_din <= x"00ac1091";
		wait for Clk_period;
		Addr <=  "0001111111111";
		Trees_din <= x"ffa41091";
		wait for Clk_period;
		Addr <=  "0010000000000";
		Trees_din <= x"08004104";
		wait for Clk_period;
		Addr <=  "0010000000001";
		Trees_din <= x"ff6a1091";
		wait for Clk_period;
		Addr <=  "0010000000010";
		Trees_din <= x"ffbd1091";
		wait for Clk_period;
		Addr <=  "0010000000011";
		Trees_din <= x"0210783c";
		wait for Clk_period;
		Addr <=  "0010000000100";
		Trees_din <= x"01fe951c";
		wait for Clk_period;
		Addr <=  "0010000000101";
		Trees_din <= x"020bce0c";
		wait for Clk_period;
		Addr <=  "0010000000110";
		Trees_din <= x"1e026a08";
		wait for Clk_period;
		Addr <=  "0010000000111";
		Trees_din <= x"1b026704";
		wait for Clk_period;
		Addr <=  "0010000001000";
		Trees_din <= x"ff821091";
		wait for Clk_period;
		Addr <=  "0010000001001";
		Trees_din <= x"008a1091";
		wait for Clk_period;
		Addr <=  "0010000001010";
		Trees_din <= x"ff551091";
		wait for Clk_period;
		Addr <=  "0010000001011";
		Trees_din <= x"0e003208";
		wait for Clk_period;
		Addr <=  "0010000001100";
		Trees_din <= x"1302ff04";
		wait for Clk_period;
		Addr <=  "0010000001101";
		Trees_din <= x"ffd31091";
		wait for Clk_period;
		Addr <=  "0010000001110";
		Trees_din <= x"009b1091";
		wait for Clk_period;
		Addr <=  "0010000001111";
		Trees_din <= x"1b027904";
		wait for Clk_period;
		Addr <=  "0010000010000";
		Trees_din <= x"ff6d1091";
		wait for Clk_period;
		Addr <=  "0010000010001";
		Trees_din <= x"00211091";
		wait for Clk_period;
		Addr <=  "0010000010010";
		Trees_din <= x"07fd1210";
		wait for Clk_period;
		Addr <=  "0010000010011";
		Trees_din <= x"0206dd08";
		wait for Clk_period;
		Addr <=  "0010000010100";
		Trees_din <= x"0d012304";
		wait for Clk_period;
		Addr <=  "0010000010101";
		Trees_din <= x"ff911091";
		wait for Clk_period;
		Addr <=  "0010000010110";
		Trees_din <= x"00261091";
		wait for Clk_period;
		Addr <=  "0010000010111";
		Trees_din <= x"0d035b04";
		wait for Clk_period;
		Addr <=  "0010000011000";
		Trees_din <= x"00191091";
		wait for Clk_period;
		Addr <=  "0010000011001";
		Trees_din <= x"ff641091";
		wait for Clk_period;
		Addr <=  "0010000011010";
		Trees_din <= x"05fb6b08";
		wait for Clk_period;
		Addr <=  "0010000011011";
		Trees_din <= x"020ab004";
		wait for Clk_period;
		Addr <=  "0010000011100";
		Trees_din <= x"00201091";
		wait for Clk_period;
		Addr <=  "0010000011101";
		Trees_din <= x"00971091";
		wait for Clk_period;
		Addr <=  "0010000011110";
		Trees_din <= x"0b007b04";
		wait for Clk_period;
		Addr <=  "0010000011111";
		Trees_din <= x"013e1091";
		wait for Clk_period;
		Addr <=  "0010000100000";
		Trees_din <= x"ffe71091";
		wait for Clk_period;
		Addr <=  "0010000100001";
		Trees_din <= x"00fd6604";
		wait for Clk_period;
		Addr <=  "0010000100010";
		Trees_din <= x"001d1091";
		wait for Clk_period;
		Addr <=  "0010000100011";
		Trees_din <= x"00971091";
		wait for Clk_period;
		Addr <=  "0010000100100";
		Trees_din <= x"01119e40";
		wait for Clk_period;
		Addr <=  "0010000100101";
		Trees_din <= x"02030518";
		wait for Clk_period;
		Addr <=  "0010000100110";
		Trees_din <= x"0800460c";
		wait for Clk_period;
		Addr <=  "0010000100111";
		Trees_din <= x"070a0704";
		wait for Clk_period;
		Addr <=  "0010000101000";
		Trees_din <= x"ff6c1115";
		wait for Clk_period;
		Addr <=  "0010000101001";
		Trees_din <= x"02017004";
		wait for Clk_period;
		Addr <=  "0010000101010";
		Trees_din <= x"ff9f1115";
		wait for Clk_period;
		Addr <=  "0010000101011";
		Trees_din <= x"00d01115";
		wait for Clk_period;
		Addr <=  "0010000101100";
		Trees_din <= x"16007408";
		wait for Clk_period;
		Addr <=  "0010000101101";
		Trees_din <= x"12008904";
		wait for Clk_period;
		Addr <=  "0010000101110";
		Trees_din <= x"012f1115";
		wait for Clk_period;
		Addr <=  "0010000101111";
		Trees_din <= x"fff61115";
		wait for Clk_period;
		Addr <=  "0010000110000";
		Trees_din <= x"ff941115";
		wait for Clk_period;
		Addr <=  "0010000110001";
		Trees_din <= x"01113d20";
		wait for Clk_period;
		Addr <=  "0010000110010";
		Trees_din <= x"02088c10";
		wait for Clk_period;
		Addr <=  "0010000110011";
		Trees_din <= x"1b024508";
		wait for Clk_period;
		Addr <=  "0010000110100";
		Trees_din <= x"01081c04";
		wait for Clk_period;
		Addr <=  "0010000110101";
		Trees_din <= x"00261115";
		wait for Clk_period;
		Addr <=  "0010000110110";
		Trees_din <= x"ff701115";
		wait for Clk_period;
		Addr <=  "0010000110111";
		Trees_din <= x"0b005a04";
		wait for Clk_period;
		Addr <=  "0010000111000";
		Trees_din <= x"00a21115";
		wait for Clk_period;
		Addr <=  "0010000111001";
		Trees_din <= x"00001115";
		wait for Clk_period;
		Addr <=  "0010000111010";
		Trees_din <= x"0d001808";
		wait for Clk_period;
		Addr <=  "0010000111011";
		Trees_din <= x"10004f04";
		wait for Clk_period;
		Addr <=  "0010000111100";
		Trees_din <= x"006a1115";
		wait for Clk_period;
		Addr <=  "0010000111101";
		Trees_din <= x"00001115";
		wait for Clk_period;
		Addr <=  "0010000111110";
		Trees_din <= x"020e3704";
		wait for Clk_period;
		Addr <=  "0010000111111";
		Trees_din <= x"000a1115";
		wait for Clk_period;
		Addr <=  "0010001000000";
		Trees_din <= x"00691115";
		wait for Clk_period;
		Addr <=  "0010001000001";
		Trees_din <= x"0b006e04";
		wait for Clk_period;
		Addr <=  "0010001000010";
		Trees_din <= x"01c11115";
		wait for Clk_period;
		Addr <=  "0010001000011";
		Trees_din <= x"ffac1115";
		wait for Clk_period;
		Addr <=  "0010001000100";
		Trees_din <= x"ff721115";
		wait for Clk_period;
		Addr <=  "0010001000101";
		Trees_din <= x"01119e28";
		wait for Clk_period;
		Addr <=  "0010001000110";
		Trees_din <= x"0200ea04";
		wait for Clk_period;
		Addr <=  "0010001000111";
		Trees_din <= x"ff781169";
		wait for Clk_period;
		Addr <=  "0010001001000";
		Trees_din <= x"1400d108";
		wait for Clk_period;
		Addr <=  "0010001001001";
		Trees_din <= x"020bce04";
		wait for Clk_period;
		Addr <=  "0010001001010";
		Trees_din <= x"ff591169";
		wait for Clk_period;
		Addr <=  "0010001001011";
		Trees_din <= x"00371169";
		wait for Clk_period;
		Addr <=  "0010001001100";
		Trees_din <= x"00117910";
		wait for Clk_period;
		Addr <=  "0010001001101";
		Trees_din <= x"1600a708";
		wait for Clk_period;
		Addr <=  "0010001001110";
		Trees_din <= x"0c008104";
		wait for Clk_period;
		Addr <=  "0010001001111";
		Trees_din <= x"004b1169";
		wait for Clk_period;
		Addr <=  "0010001010000";
		Trees_din <= x"000f1169";
		wait for Clk_period;
		Addr <=  "0010001010001";
		Trees_din <= x"07fff404";
		wait for Clk_period;
		Addr <=  "0010001010010";
		Trees_din <= x"ff6e1169";
		wait for Clk_period;
		Addr <=  "0010001010011";
		Trees_din <= x"00091169";
		wait for Clk_period;
		Addr <=  "0010001010100";
		Trees_din <= x"1401a204";
		wait for Clk_period;
		Addr <=  "0010001010101";
		Trees_din <= x"007a1169";
		wait for Clk_period;
		Addr <=  "0010001010110";
		Trees_din <= x"13040004";
		wait for Clk_period;
		Addr <=  "0010001010111";
		Trees_din <= x"ff741169";
		wait for Clk_period;
		Addr <=  "0010001011000";
		Trees_din <= x"002b1169";
		wait for Clk_period;
		Addr <=  "0010001011001";
		Trees_din <= x"ff751169";
		wait for Clk_period;
		Addr <=  "0010001011010";
		Trees_din <= x"02030518";
		wait for Clk_period;
		Addr <=  "0010001011011";
		Trees_din <= x"08004308";
		wait for Clk_period;
		Addr <=  "0010001011100";
		Trees_din <= x"01004904";
		wait for Clk_period;
		Addr <=  "0010001011101";
		Trees_din <= x"001b11dd";
		wait for Clk_period;
		Addr <=  "0010001011110";
		Trees_din <= x"ff6f11dd";
		wait for Clk_period;
		Addr <=  "0010001011111";
		Trees_din <= x"10004508";
		wait for Clk_period;
		Addr <=  "0010001100000";
		Trees_din <= x"0900b004";
		wait for Clk_period;
		Addr <=  "0010001100001";
		Trees_din <= x"000411dd";
		wait for Clk_period;
		Addr <=  "0010001100010";
		Trees_din <= x"010c11dd";
		wait for Clk_period;
		Addr <=  "0010001100011";
		Trees_din <= x"08004c04";
		wait for Clk_period;
		Addr <=  "0010001100100";
		Trees_din <= x"ff8511dd";
		wait for Clk_period;
		Addr <=  "0010001100101";
		Trees_din <= x"003e11dd";
		wait for Clk_period;
		Addr <=  "0010001100110";
		Trees_din <= x"01119e20";
		wait for Clk_period;
		Addr <=  "0010001100111";
		Trees_din <= x"0110e314";
		wait for Clk_period;
		Addr <=  "0010001101000";
		Trees_din <= x"010ff910";
		wait for Clk_period;
		Addr <=  "0010001101001";
		Trees_din <= x"0d001808";
		wait for Clk_period;
		Addr <=  "0010001101010";
		Trees_din <= x"0d000c04";
		wait for Clk_period;
		Addr <=  "0010001101011";
		Trees_din <= x"000f11dd";
		wait for Clk_period;
		Addr <=  "0010001101100";
		Trees_din <= x"005c11dd";
		wait for Clk_period;
		Addr <=  "0010001101101";
		Trees_din <= x"020a3104";
		wait for Clk_period;
		Addr <=  "0010001101110";
		Trees_din <= x"fff711dd";
		wait for Clk_period;
		Addr <=  "0010001101111";
		Trees_din <= x"002611dd";
		wait for Clk_period;
		Addr <=  "0010001110000";
		Trees_din <= x"ff7911dd";
		wait for Clk_period;
		Addr <=  "0010001110001";
		Trees_din <= x"0a004308";
		wait for Clk_period;
		Addr <=  "0010001110010";
		Trees_din <= x"05f4cf04";
		wait for Clk_period;
		Addr <=  "0010001110011";
		Trees_din <= x"006611dd";
		wait for Clk_period;
		Addr <=  "0010001110100";
		Trees_din <= x"01af11dd";
		wait for Clk_period;
		Addr <=  "0010001110101";
		Trees_din <= x"ff9811dd";
		wait for Clk_period;
		Addr <=  "0010001110110";
		Trees_din <= x"ff7e11dd";
		wait for Clk_period;
		Addr <=  "0010001110111";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0010001111000";
		Trees_din <= x"01119e44";
		wait for Clk_period;
		Addr <=  "0010001111001";
		Trees_din <= x"0200ea04";
		wait for Clk_period;
		Addr <=  "0010001111010";
		Trees_din <= x"ff7e126d";
		wait for Clk_period;
		Addr <=  "0010001111011";
		Trees_din <= x"06046d20";
		wait for Clk_period;
		Addr <=  "0010001111100";
		Trees_din <= x"020a8010";
		wait for Clk_period;
		Addr <=  "0010001111101";
		Trees_din <= x"04027f08";
		wait for Clk_period;
		Addr <=  "0010001111110";
		Trees_din <= x"03fb1b04";
		wait for Clk_period;
		Addr <=  "0010001111111";
		Trees_din <= x"001f126d";
		wait for Clk_period;
		Addr <=  "0010010000000";
		Trees_din <= x"ffe3126d";
		wait for Clk_period;
		Addr <=  "0010010000001";
		Trees_din <= x"1403f404";
		wait for Clk_period;
		Addr <=  "0010010000010";
		Trees_din <= x"000d126d";
		wait for Clk_period;
		Addr <=  "0010010000011";
		Trees_din <= x"ff7d126d";
		wait for Clk_period;
		Addr <=  "0010010000100";
		Trees_din <= x"01058308";
		wait for Clk_period;
		Addr <=  "0010010000101";
		Trees_din <= x"000b6a04";
		wait for Clk_period;
		Addr <=  "0010010000110";
		Trees_din <= x"004d126d";
		wait for Clk_period;
		Addr <=  "0010010000111";
		Trees_din <= x"ffa4126d";
		wait for Clk_period;
		Addr <=  "0010010001000";
		Trees_din <= x"0c006b04";
		wait for Clk_period;
		Addr <=  "0010010001001";
		Trees_din <= x"ff89126d";
		wait for Clk_period;
		Addr <=  "0010010001010";
		Trees_din <= x"008f126d";
		wait for Clk_period;
		Addr <=  "0010010001011";
		Trees_din <= x"1403d910";
		wait for Clk_period;
		Addr <=  "0010010001100";
		Trees_din <= x"05f3c408";
		wait for Clk_period;
		Addr <=  "0010010001101";
		Trees_din <= x"03f66c04";
		wait for Clk_period;
		Addr <=  "0010010001110";
		Trees_din <= x"ffd0126d";
		wait for Clk_period;
		Addr <=  "0010010001111";
		Trees_din <= x"0096126d";
		wait for Clk_period;
		Addr <=  "0010010010000";
		Trees_din <= x"0e003f04";
		wait for Clk_period;
		Addr <=  "0010010010001";
		Trees_din <= x"ff87126d";
		wait for Clk_period;
		Addr <=  "0010010010010";
		Trees_din <= x"0026126d";
		wait for Clk_period;
		Addr <=  "0010010010011";
		Trees_din <= x"03f84a08";
		wait for Clk_period;
		Addr <=  "0010010010100";
		Trees_din <= x"020be604";
		wait for Clk_period;
		Addr <=  "0010010010101";
		Trees_din <= x"ff9d126d";
		wait for Clk_period;
		Addr <=  "0010010010110";
		Trees_din <= x"003f126d";
		wait for Clk_period;
		Addr <=  "0010010010111";
		Trees_din <= x"01097204";
		wait for Clk_period;
		Addr <=  "0010010011000";
		Trees_din <= x"0029126d";
		wait for Clk_period;
		Addr <=  "0010010011001";
		Trees_din <= x"00e2126d";
		wait for Clk_period;
		Addr <=  "0010010011010";
		Trees_din <= x"ff7d126d";
		wait for Clk_period;
		Addr <=  "0010010011011";
		Trees_din <= x"02107868";
		wait for Clk_period;
		Addr <=  "0010010011100";
		Trees_din <= x"01fed328";
		wait for Clk_period;
		Addr <=  "0010010011101";
		Trees_din <= x"020bce14";
		wait for Clk_period;
		Addr <=  "0010010011110";
		Trees_din <= x"0e001804";
		wait for Clk_period;
		Addr <=  "0010010011111";
		Trees_din <= x"00611349";
		wait for Clk_period;
		Addr <=  "0010010100000";
		Trees_din <= x"0404c708";
		wait for Clk_period;
		Addr <=  "0010010100001";
		Trees_din <= x"020b2104";
		wait for Clk_period;
		Addr <=  "0010010100010";
		Trees_din <= x"ff5f1349";
		wait for Clk_period;
		Addr <=  "0010010100011";
		Trees_din <= x"ffe01349";
		wait for Clk_period;
		Addr <=  "0010010100100";
		Trees_din <= x"07fce404";
		wait for Clk_period;
		Addr <=  "0010010100101";
		Trees_din <= x"ffad1349";
		wait for Clk_period;
		Addr <=  "0010010100110";
		Trees_din <= x"005e1349";
		wait for Clk_period;
		Addr <=  "0010010100111";
		Trees_din <= x"0e003208";
		wait for Clk_period;
		Addr <=  "0010010101000";
		Trees_din <= x"17f84d04";
		wait for Clk_period;
		Addr <=  "0010010101001";
		Trees_din <= x"008b1349";
		wait for Clk_period;
		Addr <=  "0010010101010";
		Trees_din <= x"ffe41349";
		wait for Clk_period;
		Addr <=  "0010010101011";
		Trees_din <= x"00074808";
		wait for Clk_period;
		Addr <=  "0010010101100";
		Trees_din <= x"06085804";
		wait for Clk_period;
		Addr <=  "0010010101101";
		Trees_din <= x"00431349";
		wait for Clk_period;
		Addr <=  "0010010101110";
		Trees_din <= x"ff9d1349";
		wait for Clk_period;
		Addr <=  "0010010101111";
		Trees_din <= x"ff531349";
		wait for Clk_period;
		Addr <=  "0010010110000";
		Trees_din <= x"08003d20";
		wait for Clk_period;
		Addr <=  "0010010110001";
		Trees_din <= x"010c5210";
		wait for Clk_period;
		Addr <=  "0010010110010";
		Trees_din <= x"04067d08";
		wait for Clk_period;
		Addr <=  "0010010110011";
		Trees_din <= x"02067504";
		wait for Clk_period;
		Addr <=  "0010010110100";
		Trees_din <= x"ffc81349";
		wait for Clk_period;
		Addr <=  "0010010110101";
		Trees_din <= x"001e1349";
		wait for Clk_period;
		Addr <=  "0010010110110";
		Trees_din <= x"1b027904";
		wait for Clk_period;
		Addr <=  "0010010110111";
		Trees_din <= x"ff471349";
		wait for Clk_period;
		Addr <=  "0010010111000";
		Trees_din <= x"001f1349";
		wait for Clk_period;
		Addr <=  "0010010111001";
		Trees_din <= x"1801e508";
		wait for Clk_period;
		Addr <=  "0010010111010";
		Trees_din <= x"02094704";
		wait for Clk_period;
		Addr <=  "0010010111011";
		Trees_din <= x"ff871349";
		wait for Clk_period;
		Addr <=  "0010010111100";
		Trees_din <= x"00451349";
		wait for Clk_period;
		Addr <=  "0010010111101";
		Trees_din <= x"14034804";
		wait for Clk_period;
		Addr <=  "0010010111110";
		Trees_din <= x"ff931349";
		wait for Clk_period;
		Addr <=  "0010010111111";
		Trees_din <= x"011a1349";
		wait for Clk_period;
		Addr <=  "0010011000000";
		Trees_din <= x"15004e10";
		wait for Clk_period;
		Addr <=  "0010011000001";
		Trees_din <= x"0d000f08";
		wait for Clk_period;
		Addr <=  "0010011000010";
		Trees_din <= x"13040004";
		wait for Clk_period;
		Addr <=  "0010011000011";
		Trees_din <= x"008b1349";
		wait for Clk_period;
		Addr <=  "0010011000100";
		Trees_din <= x"00011349";
		wait for Clk_period;
		Addr <=  "0010011000101";
		Trees_din <= x"05f88f04";
		wait for Clk_period;
		Addr <=  "0010011000110";
		Trees_din <= x"00071349";
		wait for Clk_period;
		Addr <=  "0010011000111";
		Trees_din <= x"00551349";
		wait for Clk_period;
		Addr <=  "0010011001000";
		Trees_din <= x"0a004108";
		wait for Clk_period;
		Addr <=  "0010011001001";
		Trees_din <= x"07fc5704";
		wait for Clk_period;
		Addr <=  "0010011001010";
		Trees_din <= x"ffce1349";
		wait for Clk_period;
		Addr <=  "0010011001011";
		Trees_din <= x"00c31349";
		wait for Clk_period;
		Addr <=  "0010011001100";
		Trees_din <= x"18028904";
		wait for Clk_period;
		Addr <=  "0010011001101";
		Trees_din <= x"ff711349";
		wait for Clk_period;
		Addr <=  "0010011001110";
		Trees_din <= x"004b1349";
		wait for Clk_period;
		Addr <=  "0010011001111";
		Trees_din <= x"00006604";
		wait for Clk_period;
		Addr <=  "0010011010000";
		Trees_din <= x"002c1349";
		wait for Clk_period;
		Addr <=  "0010011010001";
		Trees_din <= x"00881349";
		wait for Clk_period;
		Addr <=  "0010011010010";
		Trees_din <= x"06fe0258";
		wait for Clk_period;
		Addr <=  "0010011010011";
		Trees_din <= x"1b026130";
		wait for Clk_period;
		Addr <=  "0010011010100";
		Trees_din <= x"0a004614";
		wait for Clk_period;
		Addr <=  "0010011010101";
		Trees_din <= x"0d001510";
		wait for Clk_period;
		Addr <=  "0010011010110";
		Trees_din <= x"18000d08";
		wait for Clk_period;
		Addr <=  "0010011010111";
		Trees_din <= x"04facb04";
		wait for Clk_period;
		Addr <=  "0010011011000";
		Trees_din <= x"ffe3146d";
		wait for Clk_period;
		Addr <=  "0010011011001";
		Trees_din <= x"ff74146d";
		wait for Clk_period;
		Addr <=  "0010011011010";
		Trees_din <= x"06fd5904";
		wait for Clk_period;
		Addr <=  "0010011011011";
		Trees_din <= x"ffde146d";
		wait for Clk_period;
		Addr <=  "0010011011100";
		Trees_din <= x"0084146d";
		wait for Clk_period;
		Addr <=  "0010011011101";
		Trees_din <= x"ff5e146d";
		wait for Clk_period;
		Addr <=  "0010011011110";
		Trees_din <= x"0f000510";
		wait for Clk_period;
		Addr <=  "0010011011111";
		Trees_din <= x"14040008";
		wait for Clk_period;
		Addr <=  "0010011100000";
		Trees_din <= x"01076204";
		wait for Clk_period;
		Addr <=  "0010011100001";
		Trees_din <= x"0000146d";
		wait for Clk_period;
		Addr <=  "0010011100010";
		Trees_din <= x"ff6b146d";
		wait for Clk_period;
		Addr <=  "0010011100011";
		Trees_din <= x"15003f04";
		wait for Clk_period;
		Addr <=  "0010011100100";
		Trees_din <= x"00b7146d";
		wait for Clk_period;
		Addr <=  "0010011100101";
		Trees_din <= x"ffac146d";
		wait for Clk_period;
		Addr <=  "0010011100110";
		Trees_din <= x"0b007504";
		wait for Clk_period;
		Addr <=  "0010011100111";
		Trees_din <= x"0119146d";
		wait for Clk_period;
		Addr <=  "0010011101000";
		Trees_din <= x"1100e804";
		wait for Clk_period;
		Addr <=  "0010011101001";
		Trees_din <= x"ffa5146d";
		wait for Clk_period;
		Addr <=  "0010011101010";
		Trees_din <= x"0040146d";
		wait for Clk_period;
		Addr <=  "0010011101011";
		Trees_din <= x"0704a920";
		wait for Clk_period;
		Addr <=  "0010011101100";
		Trees_din <= x"0900e910";
		wait for Clk_period;
		Addr <=  "0010011101101";
		Trees_din <= x"05f88f08";
		wait for Clk_period;
		Addr <=  "0010011101110";
		Trees_din <= x"0a005904";
		wait for Clk_period;
		Addr <=  "0010011101111";
		Trees_din <= x"0001146d";
		wait for Clk_period;
		Addr <=  "0010011110000";
		Trees_din <= x"00e9146d";
		wait for Clk_period;
		Addr <=  "0010011110001";
		Trees_din <= x"01fbed04";
		wait for Clk_period;
		Addr <=  "0010011110010";
		Trees_din <= x"ffd0146d";
		wait for Clk_period;
		Addr <=  "0010011110011";
		Trees_din <= x"00bc146d";
		wait for Clk_period;
		Addr <=  "0010011110100";
		Trees_din <= x"0e002508";
		wait for Clk_period;
		Addr <=  "0010011110101";
		Trees_din <= x"18000d04";
		wait for Clk_period;
		Addr <=  "0010011110110";
		Trees_din <= x"0031146d";
		wait for Clk_period;
		Addr <=  "0010011110111";
		Trees_din <= x"ff94146d";
		wait for Clk_period;
		Addr <=  "0010011111000";
		Trees_din <= x"0a004004";
		wait for Clk_period;
		Addr <=  "0010011111001";
		Trees_din <= x"0034146d";
		wait for Clk_period;
		Addr <=  "0010011111010";
		Trees_din <= x"0160146d";
		wait for Clk_period;
		Addr <=  "0010011111011";
		Trees_din <= x"0a003e04";
		wait for Clk_period;
		Addr <=  "0010011111100";
		Trees_din <= x"0030146d";
		wait for Clk_period;
		Addr <=  "0010011111101";
		Trees_din <= x"ff72146d";
		wait for Clk_period;
		Addr <=  "0010011111110";
		Trees_din <= x"03fc4020";
		wait for Clk_period;
		Addr <=  "0010011111111";
		Trees_din <= x"08004d14";
		wait for Clk_period;
		Addr <=  "0010100000000";
		Trees_din <= x"02024504";
		wait for Clk_period;
		Addr <=  "0010100000001";
		Trees_din <= x"ff7c146d";
		wait for Clk_period;
		Addr <=  "0010100000010";
		Trees_din <= x"04fdcc08";
		wait for Clk_period;
		Addr <=  "0010100000011";
		Trees_din <= x"04fc6804";
		wait for Clk_period;
		Addr <=  "0010100000100";
		Trees_din <= x"ffe8146d";
		wait for Clk_period;
		Addr <=  "0010100000101";
		Trees_din <= x"0061146d";
		wait for Clk_period;
		Addr <=  "0010100000110";
		Trees_din <= x"010dfe04";
		wait for Clk_period;
		Addr <=  "0010100000111";
		Trees_din <= x"0004146d";
		wait for Clk_period;
		Addr <=  "0010100001000";
		Trees_din <= x"ffa3146d";
		wait for Clk_period;
		Addr <=  "0010100001001";
		Trees_din <= x"1c028708";
		wait for Clk_period;
		Addr <=  "0010100001010";
		Trees_din <= x"15004a04";
		wait for Clk_period;
		Addr <=  "0010100001011";
		Trees_din <= x"ff46146d";
		wait for Clk_period;
		Addr <=  "0010100001100";
		Trees_din <= x"ffd6146d";
		wait for Clk_period;
		Addr <=  "0010100001101";
		Trees_din <= x"0035146d";
		wait for Clk_period;
		Addr <=  "0010100001110";
		Trees_din <= x"02097f14";
		wait for Clk_period;
		Addr <=  "0010100001111";
		Trees_din <= x"20040008";
		wait for Clk_period;
		Addr <=  "0010100010000";
		Trees_din <= x"03fe6004";
		wait for Clk_period;
		Addr <=  "0010100010001";
		Trees_din <= x"fffb146d";
		wait for Clk_period;
		Addr <=  "0010100010010";
		Trees_din <= x"0070146d";
		wait for Clk_period;
		Addr <=  "0010100010011";
		Trees_din <= x"00006604";
		wait for Clk_period;
		Addr <=  "0010100010100";
		Trees_din <= x"0004146d";
		wait for Clk_period;
		Addr <=  "0010100010101";
		Trees_din <= x"19000a04";
		wait for Clk_period;
		Addr <=  "0010100010110";
		Trees_din <= x"ff3a146d";
		wait for Clk_period;
		Addr <=  "0010100010111";
		Trees_din <= x"ffd8146d";
		wait for Clk_period;
		Addr <=  "0010100011000";
		Trees_din <= x"01010e04";
		wait for Clk_period;
		Addr <=  "0010100011001";
		Trees_din <= x"ffc7146d";
		wait for Clk_period;
		Addr <=  "0010100011010";
		Trees_din <= x"0086146d";
		wait for Clk_period;
		Addr <=  "0010100011011";
		Trees_din <= x"02107864";
		wait for Clk_period;
		Addr <=  "0010100011100";
		Trees_din <= x"06046d40";
		wait for Clk_period;
		Addr <=  "0010100011101";
		Trees_din <= x"02088c20";
		wait for Clk_period;
		Addr <=  "0010100011110";
		Trees_din <= x"08003a10";
		wait for Clk_period;
		Addr <=  "0010100011111";
		Trees_din <= x"1d028008";
		wait for Clk_period;
		Addr <=  "0010100100000";
		Trees_din <= x"10005604";
		wait for Clk_period;
		Addr <=  "0010100100001";
		Trees_din <= x"ff9f1541";
		wait for Clk_period;
		Addr <=  "0010100100010";
		Trees_din <= x"00311541";
		wait for Clk_period;
		Addr <=  "0010100100011";
		Trees_din <= x"06ffff04";
		wait for Clk_period;
		Addr <=  "0010100100100";
		Trees_din <= x"008d1541";
		wait for Clk_period;
		Addr <=  "0010100100101";
		Trees_din <= x"ff7d1541";
		wait for Clk_period;
		Addr <=  "0010100100110";
		Trees_din <= x"000bff08";
		wait for Clk_period;
		Addr <=  "0010100100111";
		Trees_din <= x"03f63104";
		wait for Clk_period;
		Addr <=  "0010100101000";
		Trees_din <= x"00a91541";
		wait for Clk_period;
		Addr <=  "0010100101001";
		Trees_din <= x"000d1541";
		wait for Clk_period;
		Addr <=  "0010100101010";
		Trees_din <= x"10003f04";
		wait for Clk_period;
		Addr <=  "0010100101011";
		Trees_din <= x"004b1541";
		wait for Clk_period;
		Addr <=  "0010100101100";
		Trees_din <= x"ffa41541";
		wait for Clk_period;
		Addr <=  "0010100101101";
		Trees_din <= x"04025f10";
		wait for Clk_period;
		Addr <=  "0010100101110";
		Trees_din <= x"15004e08";
		wait for Clk_period;
		Addr <=  "0010100101111";
		Trees_din <= x"11006404";
		wait for Clk_period;
		Addr <=  "0010100110000";
		Trees_din <= x"00941541";
		wait for Clk_period;
		Addr <=  "0010100110001";
		Trees_din <= x"00251541";
		wait for Clk_period;
		Addr <=  "0010100110010";
		Trees_din <= x"07ff7e04";
		wait for Clk_period;
		Addr <=  "0010100110011";
		Trees_din <= x"ff7a1541";
		wait for Clk_period;
		Addr <=  "0010100110100";
		Trees_din <= x"005a1541";
		wait for Clk_period;
		Addr <=  "0010100110101";
		Trees_din <= x"0a003c08";
		wait for Clk_period;
		Addr <=  "0010100110110";
		Trees_din <= x"08003f04";
		wait for Clk_period;
		Addr <=  "0010100110111";
		Trees_din <= x"ffde1541";
		wait for Clk_period;
		Addr <=  "0010100111000";
		Trees_din <= x"00b91541";
		wait for Clk_period;
		Addr <=  "0010100111001";
		Trees_din <= x"17f7c004";
		wait for Clk_period;
		Addr <=  "0010100111010";
		Trees_din <= x"ffa31541";
		wait for Clk_period;
		Addr <=  "0010100111011";
		Trees_din <= x"00041541";
		wait for Clk_period;
		Addr <=  "0010100111100";
		Trees_din <= x"03fb421c";
		wait for Clk_period;
		Addr <=  "0010100111101";
		Trees_din <= x"1000440c";
		wait for Clk_period;
		Addr <=  "0010100111110";
		Trees_din <= x"16006408";
		wait for Clk_period;
		Addr <=  "0010100111111";
		Trees_din <= x"1f027c04";
		wait for Clk_period;
		Addr <=  "0010101000000";
		Trees_din <= x"000b1541";
		wait for Clk_period;
		Addr <=  "0010101000001";
		Trees_din <= x"ff7b1541";
		wait for Clk_period;
		Addr <=  "0010101000010";
		Trees_din <= x"ff321541";
		wait for Clk_period;
		Addr <=  "0010101000011";
		Trees_din <= x"00071e08";
		wait for Clk_period;
		Addr <=  "0010101000100";
		Trees_din <= x"0206c404";
		wait for Clk_period;
		Addr <=  "0010101000101";
		Trees_din <= x"ff801541";
		wait for Clk_period;
		Addr <=  "0010101000110";
		Trees_din <= x"00301541";
		wait for Clk_period;
		Addr <=  "0010101000111";
		Trees_din <= x"020bce04";
		wait for Clk_period;
		Addr <=  "0010101001000";
		Trees_din <= x"ff7b1541";
		wait for Clk_period;
		Addr <=  "0010101001001";
		Trees_din <= x"000d1541";
		wait for Clk_period;
		Addr <=  "0010101001010";
		Trees_din <= x"10003f04";
		wait for Clk_period;
		Addr <=  "0010101001011";
		Trees_din <= x"00041541";
		wait for Clk_period;
		Addr <=  "0010101001100";
		Trees_din <= x"00c71541";
		wait for Clk_period;
		Addr <=  "0010101001101";
		Trees_din <= x"17f77a04";
		wait for Clk_period;
		Addr <=  "0010101001110";
		Trees_din <= x"00241541";
		wait for Clk_period;
		Addr <=  "0010101001111";
		Trees_din <= x"00831541";
		wait for Clk_period;
		Addr <=  "0010101010000";
		Trees_din <= x"1400d108";
		wait for Clk_period;
		Addr <=  "0010101010001";
		Trees_din <= x"020bce04";
		wait for Clk_period;
		Addr <=  "0010101010010";
		Trees_din <= x"ff66163d";
		wait for Clk_period;
		Addr <=  "0010101010011";
		Trees_din <= x"0031163d";
		wait for Clk_period;
		Addr <=  "0010101010100";
		Trees_din <= x"06fe0240";
		wait for Clk_period;
		Addr <=  "0010101010101";
		Trees_din <= x"1e025f20";
		wait for Clk_period;
		Addr <=  "0010101010110";
		Trees_din <= x"06fd3710";
		wait for Clk_period;
		Addr <=  "0010101010111";
		Trees_din <= x"0a004808";
		wait for Clk_period;
		Addr <=  "0010101011000";
		Trees_din <= x"02096b04";
		wait for Clk_period;
		Addr <=  "0010101011001";
		Trees_din <= x"ff65163d";
		wait for Clk_period;
		Addr <=  "0010101011010";
		Trees_din <= x"ffeb163d";
		wait for Clk_period;
		Addr <=  "0010101011011";
		Trees_din <= x"0c00a804";
		wait for Clk_period;
		Addr <=  "0010101011100";
		Trees_din <= x"ffba163d";
		wait for Clk_period;
		Addr <=  "0010101011101";
		Trees_din <= x"005d163d";
		wait for Clk_period;
		Addr <=  "0010101011110";
		Trees_din <= x"15003e08";
		wait for Clk_period;
		Addr <=  "0010101011111";
		Trees_din <= x"0d000604";
		wait for Clk_period;
		Addr <=  "0010101100000";
		Trees_din <= x"0033163d";
		wait for Clk_period;
		Addr <=  "0010101100001";
		Trees_din <= x"ff73163d";
		wait for Clk_period;
		Addr <=  "0010101100010";
		Trees_din <= x"15003f04";
		wait for Clk_period;
		Addr <=  "0010101100011";
		Trees_din <= x"015c163d";
		wait for Clk_period;
		Addr <=  "0010101100100";
		Trees_din <= x"0021163d";
		wait for Clk_period;
		Addr <=  "0010101100101";
		Trees_din <= x"1c027210";
		wait for Clk_period;
		Addr <=  "0010101100110";
		Trees_din <= x"04fdd608";
		wait for Clk_period;
		Addr <=  "0010101100111";
		Trees_din <= x"06fdde04";
		wait for Clk_period;
		Addr <=  "0010101101000";
		Trees_din <= x"0004163d";
		wait for Clk_period;
		Addr <=  "0010101101001";
		Trees_din <= x"0147163d";
		wait for Clk_period;
		Addr <=  "0010101101010";
		Trees_din <= x"0c00ae04";
		wait for Clk_period;
		Addr <=  "0010101101011";
		Trees_din <= x"00ef163d";
		wait for Clk_period;
		Addr <=  "0010101101100";
		Trees_din <= x"000f163d";
		wait for Clk_period;
		Addr <=  "0010101101101";
		Trees_din <= x"05f82f08";
		wait for Clk_period;
		Addr <=  "0010101101110";
		Trees_din <= x"19001904";
		wait for Clk_period;
		Addr <=  "0010101101111";
		Trees_din <= x"ffb7163d";
		wait for Clk_period;
		Addr <=  "0010101110000";
		Trees_din <= x"0070163d";
		wait for Clk_period;
		Addr <=  "0010101110001";
		Trees_din <= x"0d007004";
		wait for Clk_period;
		Addr <=  "0010101110010";
		Trees_din <= x"ffc9163d";
		wait for Clk_period;
		Addr <=  "0010101110011";
		Trees_din <= x"009a163d";
		wait for Clk_period;
		Addr <=  "0010101110100";
		Trees_din <= x"0d00011c";
		wait for Clk_period;
		Addr <=  "0010101110101";
		Trees_din <= x"1f024d0c";
		wait for Clk_period;
		Addr <=  "0010101110110";
		Trees_din <= x"0209bd04";
		wait for Clk_period;
		Addr <=  "0010101110111";
		Trees_din <= x"ff5b163d";
		wait for Clk_period;
		Addr <=  "0010101111000";
		Trees_din <= x"1b024804";
		wait for Clk_period;
		Addr <=  "0010101111001";
		Trees_din <= x"0075163d";
		wait for Clk_period;
		Addr <=  "0010101111010";
		Trees_din <= x"ffe5163d";
		wait for Clk_period;
		Addr <=  "0010101111011";
		Trees_din <= x"010c9108";
		wait for Clk_period;
		Addr <=  "0010101111100";
		Trees_din <= x"03f74904";
		wait for Clk_period;
		Addr <=  "0010101111101";
		Trees_din <= x"ffef163d";
		wait for Clk_period;
		Addr <=  "0010101111110";
		Trees_din <= x"00ba163d";
		wait for Clk_period;
		Addr <=  "0010101111111";
		Trees_din <= x"1403fd04";
		wait for Clk_period;
		Addr <=  "0010110000000";
		Trees_din <= x"0028163d";
		wait for Clk_period;
		Addr <=  "0010110000001";
		Trees_din <= x"ff8d163d";
		wait for Clk_period;
		Addr <=  "0010110000010";
		Trees_din <= x"03fc4010";
		wait for Clk_period;
		Addr <=  "0010110000011";
		Trees_din <= x"0900e108";
		wait for Clk_period;
		Addr <=  "0010110000100";
		Trees_din <= x"0900c004";
		wait for Clk_period;
		Addr <=  "0010110000101";
		Trees_din <= x"fff4163d";
		wait for Clk_period;
		Addr <=  "0010110000110";
		Trees_din <= x"0030163d";
		wait for Clk_period;
		Addr <=  "0010110000111";
		Trees_din <= x"07f81804";
		wait for Clk_period;
		Addr <=  "0010110001000";
		Trees_din <= x"0058163d";
		wait for Clk_period;
		Addr <=  "0010110001001";
		Trees_din <= x"ffc9163d";
		wait for Clk_period;
		Addr <=  "0010110001010";
		Trees_din <= x"20040004";
		wait for Clk_period;
		Addr <=  "0010110001011";
		Trees_din <= x"0047163d";
		wait for Clk_period;
		Addr <=  "0010110001100";
		Trees_din <= x"02097f04";
		wait for Clk_period;
		Addr <=  "0010110001101";
		Trees_din <= x"ff59163d";
		wait for Clk_period;
		Addr <=  "0010110001110";
		Trees_din <= x"002c163d";
		wait for Clk_period;
		Addr <=  "0010110001111";
		Trees_din <= x"1ff9b004";
		wait for Clk_period;
		Addr <=  "0010110010000";
		Trees_din <= x"ff821709";
		wait for Clk_period;
		Addr <=  "0010110010001";
		Trees_din <= x"12008640";
		wait for Clk_period;
		Addr <=  "0010110010010";
		Trees_din <= x"0204ff20";
		wait for Clk_period;
		Addr <=  "0010110010011";
		Trees_din <= x"05f8d210";
		wait for Clk_period;
		Addr <=  "0010110010100";
		Trees_din <= x"0900e908";
		wait for Clk_period;
		Addr <=  "0010110010101";
		Trees_din <= x"1af94c04";
		wait for Clk_period;
		Addr <=  "0010110010110";
		Trees_din <= x"00251709";
		wait for Clk_period;
		Addr <=  "0010110010111";
		Trees_din <= x"ff7e1709";
		wait for Clk_period;
		Addr <=  "0010110011000";
		Trees_din <= x"0203b504";
		wait for Clk_period;
		Addr <=  "0010110011001";
		Trees_din <= x"ff8d1709";
		wait for Clk_period;
		Addr <=  "0010110011010";
		Trees_din <= x"006a1709";
		wait for Clk_period;
		Addr <=  "0010110011011";
		Trees_din <= x"1afc5408";
		wait for Clk_period;
		Addr <=  "0010110011100";
		Trees_din <= x"05fad604";
		wait for Clk_period;
		Addr <=  "0010110011101";
		Trees_din <= x"00a71709";
		wait for Clk_period;
		Addr <=  "0010110011110";
		Trees_din <= x"ffe31709";
		wait for Clk_period;
		Addr <=  "0010110011111";
		Trees_din <= x"01008904";
		wait for Clk_period;
		Addr <=  "0010110100000";
		Trees_din <= x"fff21709";
		wait for Clk_period;
		Addr <=  "0010110100001";
		Trees_din <= x"ff7f1709";
		wait for Clk_period;
		Addr <=  "0010110100010";
		Trees_din <= x"10004410";
		wait for Clk_period;
		Addr <=  "0010110100011";
		Trees_din <= x"0900b508";
		wait for Clk_period;
		Addr <=  "0010110100100";
		Trees_din <= x"0d000704";
		wait for Clk_period;
		Addr <=  "0010110100101";
		Trees_din <= x"00241709";
		wait for Clk_period;
		Addr <=  "0010110100110";
		Trees_din <= x"ff431709";
		wait for Clk_period;
		Addr <=  "0010110100111";
		Trees_din <= x"17f70f04";
		wait for Clk_period;
		Addr <=  "0010110101000";
		Trees_din <= x"007d1709";
		wait for Clk_period;
		Addr <=  "0010110101001";
		Trees_din <= x"ffec1709";
		wait for Clk_period;
		Addr <=  "0010110101010";
		Trees_din <= x"10004808";
		wait for Clk_period;
		Addr <=  "0010110101011";
		Trees_din <= x"1302e704";
		wait for Clk_period;
		Addr <=  "0010110101100";
		Trees_din <= x"ffd51709";
		wait for Clk_period;
		Addr <=  "0010110101101";
		Trees_din <= x"006a1709";
		wait for Clk_period;
		Addr <=  "0010110101110";
		Trees_din <= x"12008204";
		wait for Clk_period;
		Addr <=  "0010110101111";
		Trees_din <= x"00101709";
		wait for Clk_period;
		Addr <=  "0010110110000";
		Trees_din <= x"ff921709";
		wait for Clk_period;
		Addr <=  "0010110110001";
		Trees_din <= x"1af9c10c";
		wait for Clk_period;
		Addr <=  "0010110110010";
		Trees_din <= x"06fd1a04";
		wait for Clk_period;
		Addr <=  "0010110110011";
		Trees_din <= x"00291709";
		wait for Clk_period;
		Addr <=  "0010110110100";
		Trees_din <= x"01039604";
		wait for Clk_period;
		Addr <=  "0010110110101";
		Trees_din <= x"ffe51709";
		wait for Clk_period;
		Addr <=  "0010110110110";
		Trees_din <= x"ff5d1709";
		wait for Clk_period;
		Addr <=  "0010110110111";
		Trees_din <= x"13039a0c";
		wait for Clk_period;
		Addr <=  "0010110111000";
		Trees_din <= x"0e003408";
		wait for Clk_period;
		Addr <=  "0010110111001";
		Trees_din <= x"0d035b04";
		wait for Clk_period;
		Addr <=  "0010110111010";
		Trees_din <= x"008c1709";
		wait for Clk_period;
		Addr <=  "0010110111011";
		Trees_din <= x"ffdb1709";
		wait for Clk_period;
		Addr <=  "0010110111100";
		Trees_din <= x"ff7a1709";
		wait for Clk_period;
		Addr <=  "0010110111101";
		Trees_din <= x"07f97504";
		wait for Clk_period;
		Addr <=  "0010110111110";
		Trees_din <= x"ff661709";
		wait for Clk_period;
		Addr <=  "0010110111111";
		Trees_din <= x"02079a04";
		wait for Clk_period;
		Addr <=  "0010111000000";
		Trees_din <= x"ffe71709";
		wait for Clk_period;
		Addr <=  "0010111000001";
		Trees_din <= x"006f1709";
		wait for Clk_period;
		Addr <=  "0010111000010";
		Trees_din <= x"0600b778";
		wait for Clk_period;
		Addr <=  "0010111000011";
		Trees_din <= x"08003e40";
		wait for Clk_period;
		Addr <=  "0010111000100";
		Trees_din <= x"0207f120";
		wait for Clk_period;
		Addr <=  "0010111000101";
		Trees_din <= x"1b028010";
		wait for Clk_period;
		Addr <=  "0010111000110";
		Trees_din <= x"05f72708";
		wait for Clk_period;
		Addr <=  "0010111000111";
		Trees_din <= x"08003004";
		wait for Clk_period;
		Addr <=  "0010111001000";
		Trees_din <= x"ffee189d";
		wait for Clk_period;
		Addr <=  "0010111001001";
		Trees_din <= x"ff7f189d";
		wait for Clk_period;
		Addr <=  "0010111001010";
		Trees_din <= x"0205ec04";
		wait for Clk_period;
		Addr <=  "0010111001011";
		Trees_din <= x"ff95189d";
		wait for Clk_period;
		Addr <=  "0010111001100";
		Trees_din <= x"004e189d";
		wait for Clk_period;
		Addr <=  "0010111001101";
		Trees_din <= x"0700f908";
		wait for Clk_period;
		Addr <=  "0010111001110";
		Trees_din <= x"0b008f04";
		wait for Clk_period;
		Addr <=  "0010111001111";
		Trees_din <= x"0083189d";
		wait for Clk_period;
		Addr <=  "0010111010000";
		Trees_din <= x"ffcc189d";
		wait for Clk_period;
		Addr <=  "0010111010001";
		Trees_din <= x"03fc5c04";
		wait for Clk_period;
		Addr <=  "0010111010010";
		Trees_din <= x"ff90189d";
		wait for Clk_period;
		Addr <=  "0010111010011";
		Trees_din <= x"ffe1189d";
		wait for Clk_period;
		Addr <=  "0010111010100";
		Trees_din <= x"05f5f610";
		wait for Clk_period;
		Addr <=  "0010111010101";
		Trees_din <= x"07ff6f08";
		wait for Clk_period;
		Addr <=  "0010111010110";
		Trees_din <= x"01095e04";
		wait for Clk_period;
		Addr <=  "0010111010111";
		Trees_din <= x"ff57189d";
		wait for Clk_period;
		Addr <=  "0010111011000";
		Trees_din <= x"fff9189d";
		wait for Clk_period;
		Addr <=  "0010111011001";
		Trees_din <= x"1f024b04";
		wait for Clk_period;
		Addr <=  "0010111011010";
		Trees_din <= x"000b189d";
		wait for Clk_period;
		Addr <=  "0010111011011";
		Trees_din <= x"0086189d";
		wait for Clk_period;
		Addr <=  "0010111011100";
		Trees_din <= x"03fc1e08";
		wait for Clk_period;
		Addr <=  "0010111011101";
		Trees_din <= x"04007504";
		wait for Clk_period;
		Addr <=  "0010111011110";
		Trees_din <= x"00db189d";
		wait for Clk_period;
		Addr <=  "0010111011111";
		Trees_din <= x"0026189d";
		wait for Clk_period;
		Addr <=  "0010111100000";
		Trees_din <= x"10004404";
		wait for Clk_period;
		Addr <=  "0010111100001";
		Trees_din <= x"ff91189d";
		wait for Clk_period;
		Addr <=  "0010111100010";
		Trees_din <= x"006f189d";
		wait for Clk_period;
		Addr <=  "0010111100011";
		Trees_din <= x"0a00421c";
		wait for Clk_period;
		Addr <=  "0010111100100";
		Trees_din <= x"0900bf0c";
		wait for Clk_period;
		Addr <=  "0010111100101";
		Trees_din <= x"0a003e08";
		wait for Clk_period;
		Addr <=  "0010111100110";
		Trees_din <= x"0a003e04";
		wait for Clk_period;
		Addr <=  "0010111100111";
		Trees_din <= x"ffaf189d";
		wait for Clk_period;
		Addr <=  "0010111101000";
		Trees_din <= x"0090189d";
		wait for Clk_period;
		Addr <=  "0010111101001";
		Trees_din <= x"ff71189d";
		wait for Clk_period;
		Addr <=  "0010111101010";
		Trees_din <= x"0900dc08";
		wait for Clk_period;
		Addr <=  "0010111101011";
		Trees_din <= x"0a003f04";
		wait for Clk_period;
		Addr <=  "0010111101100";
		Trees_din <= x"0009189d";
		wait for Clk_period;
		Addr <=  "0010111101101";
		Trees_din <= x"0134189d";
		wait for Clk_period;
		Addr <=  "0010111101110";
		Trees_din <= x"08004504";
		wait for Clk_period;
		Addr <=  "0010111101111";
		Trees_din <= x"0049189d";
		wait for Clk_period;
		Addr <=  "0010111110000";
		Trees_din <= x"ff7a189d";
		wait for Clk_period;
		Addr <=  "0010111110001";
		Trees_din <= x"0b00670c";
		wait for Clk_period;
		Addr <=  "0010111110010";
		Trees_din <= x"08004c08";
		wait for Clk_period;
		Addr <=  "0010111110011";
		Trees_din <= x"0c006e04";
		wait for Clk_period;
		Addr <=  "0010111110100";
		Trees_din <= x"0019189d";
		wait for Clk_period;
		Addr <=  "0010111110101";
		Trees_din <= x"ff5e189d";
		wait for Clk_period;
		Addr <=  "0010111110110";
		Trees_din <= x"005c189d";
		wait for Clk_period;
		Addr <=  "0010111110111";
		Trees_din <= x"1b027a08";
		wait for Clk_period;
		Addr <=  "0010111111000";
		Trees_din <= x"01093504";
		wait for Clk_period;
		Addr <=  "0010111111001";
		Trees_din <= x"fff8189d";
		wait for Clk_period;
		Addr <=  "0010111111010";
		Trees_din <= x"0072189d";
		wait for Clk_period;
		Addr <=  "0010111111011";
		Trees_din <= x"06fbf104";
		wait for Clk_period;
		Addr <=  "0010111111100";
		Trees_din <= x"0030189d";
		wait for Clk_period;
		Addr <=  "0010111111101";
		Trees_din <= x"ffa6189d";
		wait for Clk_period;
		Addr <=  "0010111111110";
		Trees_din <= x"0d000120";
		wait for Clk_period;
		Addr <=  "0010111111111";
		Trees_din <= x"1b02560c";
		wait for Clk_period;
		Addr <=  "0011000000000";
		Trees_din <= x"1d023004";
		wait for Clk_period;
		Addr <=  "0011000000001";
		Trees_din <= x"0021189d";
		wait for Clk_period;
		Addr <=  "0011000000010";
		Trees_din <= x"1afd5e04";
		wait for Clk_period;
		Addr <=  "0011000000011";
		Trees_din <= x"fff3189d";
		wait for Clk_period;
		Addr <=  "0011000000100";
		Trees_din <= x"ff7f189d";
		wait for Clk_period;
		Addr <=  "0011000000101";
		Trees_din <= x"0c00ab0c";
		wait for Clk_period;
		Addr <=  "0011000000110";
		Trees_din <= x"03f82708";
		wait for Clk_period;
		Addr <=  "0011000000111";
		Trees_din <= x"07f79c04";
		wait for Clk_period;
		Addr <=  "0011000001000";
		Trees_din <= x"00ac189d";
		wait for Clk_period;
		Addr <=  "0011000001001";
		Trees_din <= x"fff9189d";
		wait for Clk_period;
		Addr <=  "0011000001010";
		Trees_din <= x"00d4189d";
		wait for Clk_period;
		Addr <=  "0011000001011";
		Trees_din <= x"19000f04";
		wait for Clk_period;
		Addr <=  "0011000001100";
		Trees_din <= x"ffe6189d";
		wait for Clk_period;
		Addr <=  "0011000001101";
		Trees_din <= x"0037189d";
		wait for Clk_period;
		Addr <=  "0011000001110";
		Trees_din <= x"06011914";
		wait for Clk_period;
		Addr <=  "0011000001111";
		Trees_din <= x"010f6410";
		wait for Clk_period;
		Addr <=  "0011000010000";
		Trees_din <= x"0403b208";
		wait for Clk_period;
		Addr <=  "0011000010001";
		Trees_din <= x"05f86604";
		wait for Clk_period;
		Addr <=  "0011000010010";
		Trees_din <= x"ff49189d";
		wait for Clk_period;
		Addr <=  "0011000010011";
		Trees_din <= x"ffe4189d";
		wait for Clk_period;
		Addr <=  "0011000010100";
		Trees_din <= x"03f7e704";
		wait for Clk_period;
		Addr <=  "0011000010101";
		Trees_din <= x"ffaa189d";
		wait for Clk_period;
		Addr <=  "0011000010110";
		Trees_din <= x"006d189d";
		wait for Clk_period;
		Addr <=  "0011000010111";
		Trees_din <= x"009a189d";
		wait for Clk_period;
		Addr <=  "0011000011000";
		Trees_din <= x"05f3e610";
		wait for Clk_period;
		Addr <=  "0011000011001";
		Trees_din <= x"010ca908";
		wait for Clk_period;
		Addr <=  "0011000011010";
		Trees_din <= x"0900e404";
		wait for Clk_period;
		Addr <=  "0011000011011";
		Trees_din <= x"0085189d";
		wait for Clk_period;
		Addr <=  "0011000011100";
		Trees_din <= x"ffca189d";
		wait for Clk_period;
		Addr <=  "0011000011101";
		Trees_din <= x"0b008204";
		wait for Clk_period;
		Addr <=  "0011000011110";
		Trees_din <= x"ff72189d";
		wait for Clk_period;
		Addr <=  "0011000011111";
		Trees_din <= x"002b189d";
		wait for Clk_period;
		Addr <=  "0011000100000";
		Trees_din <= x"05f58408";
		wait for Clk_period;
		Addr <=  "0011000100001";
		Trees_din <= x"03f8d704";
		wait for Clk_period;
		Addr <=  "0011000100010";
		Trees_din <= x"ff7c189d";
		wait for Clk_period;
		Addr <=  "0011000100011";
		Trees_din <= x"0008189d";
		wait for Clk_period;
		Addr <=  "0011000100100";
		Trees_din <= x"0a003f04";
		wait for Clk_period;
		Addr <=  "0011000100101";
		Trees_din <= x"0030189d";
		wait for Clk_period;
		Addr <=  "0011000100110";
		Trees_din <= x"ffee189d";
		wait for Clk_period;
		Addr <=  "0011000100111";
		Trees_din <= x"0210786c";
		wait for Clk_period;
		Addr <=  "0011000101000";
		Trees_din <= x"0600c038";
		wait for Clk_period;
		Addr <=  "0011000101001";
		Trees_din <= x"0a00501c";
		wait for Clk_period;
		Addr <=  "0011000101010";
		Trees_din <= x"03fb1b0c";
		wait for Clk_period;
		Addr <=  "0011000101011";
		Trees_din <= x"07057108";
		wait for Clk_period;
		Addr <=  "0011000101100";
		Trees_din <= x"0400d004";
		wait for Clk_period;
		Addr <=  "0011000101101";
		Trees_din <= x"003a1981";
		wait for Clk_period;
		Addr <=  "0011000101110";
		Trees_din <= x"fff81981";
		wait for Clk_period;
		Addr <=  "0011000101111";
		Trees_din <= x"ff7e1981";
		wait for Clk_period;
		Addr <=  "0011000110000";
		Trees_din <= x"0900a908";
		wait for Clk_period;
		Addr <=  "0011000110001";
		Trees_din <= x"1f027604";
		wait for Clk_period;
		Addr <=  "0011000110010";
		Trees_din <= x"00761981";
		wait for Clk_period;
		Addr <=  "0011000110011";
		Trees_din <= x"ffda1981";
		wait for Clk_period;
		Addr <=  "0011000110100";
		Trees_din <= x"04f77004";
		wait for Clk_period;
		Addr <=  "0011000110101";
		Trees_din <= x"005c1981";
		wait for Clk_period;
		Addr <=  "0011000110110";
		Trees_din <= x"ffb71981";
		wait for Clk_period;
		Addr <=  "0011000110111";
		Trees_din <= x"0a005910";
		wait for Clk_period;
		Addr <=  "0011000111000";
		Trees_din <= x"0105e908";
		wait for Clk_period;
		Addr <=  "0011000111001";
		Trees_din <= x"08003e04";
		wait for Clk_period;
		Addr <=  "0011000111010";
		Trees_din <= x"004c1981";
		wait for Clk_period;
		Addr <=  "0011000111011";
		Trees_din <= x"ffe01981";
		wait for Clk_period;
		Addr <=  "0011000111100";
		Trees_din <= x"1b048204";
		wait for Clk_period;
		Addr <=  "0011000111101";
		Trees_din <= x"ff761981";
		wait for Clk_period;
		Addr <=  "0011000111110";
		Trees_din <= x"00171981";
		wait for Clk_period;
		Addr <=  "0011000111111";
		Trees_din <= x"0b008404";
		wait for Clk_period;
		Addr <=  "0011001000000";
		Trees_din <= x"00bc1981";
		wait for Clk_period;
		Addr <=  "0011001000001";
		Trees_din <= x"01081c04";
		wait for Clk_period;
		Addr <=  "0011001000010";
		Trees_din <= x"00041981";
		wait for Clk_period;
		Addr <=  "0011001000011";
		Trees_din <= x"ff8a1981";
		wait for Clk_period;
		Addr <=  "0011001000100";
		Trees_din <= x"06011914";
		wait for Clk_period;
		Addr <=  "0011001000101";
		Trees_din <= x"020a310c";
		wait for Clk_period;
		Addr <=  "0011001000110";
		Trees_din <= x"010f7d08";
		wait for Clk_period;
		Addr <=  "0011001000111";
		Trees_din <= x"01076204";
		wait for Clk_period;
		Addr <=  "0011001001000";
		Trees_din <= x"fff01981";
		wait for Clk_period;
		Addr <=  "0011001001001";
		Trees_din <= x"ff5b1981";
		wait for Clk_period;
		Addr <=  "0011001001010";
		Trees_din <= x"001d1981";
		wait for Clk_period;
		Addr <=  "0011001001011";
		Trees_din <= x"08003e04";
		wait for Clk_period;
		Addr <=  "0011001001100";
		Trees_din <= x"ffc01981";
		wait for Clk_period;
		Addr <=  "0011001001101";
		Trees_din <= x"006f1981";
		wait for Clk_period;
		Addr <=  "0011001001110";
		Trees_din <= x"03f92810";
		wait for Clk_period;
		Addr <=  "0011001001111";
		Trees_din <= x"0208b708";
		wait for Clk_period;
		Addr <=  "0011001010000";
		Trees_din <= x"07fbfd04";
		wait for Clk_period;
		Addr <=  "0011001010001";
		Trees_din <= x"ff691981";
		wait for Clk_period;
		Addr <=  "0011001010010";
		Trees_din <= x"ffee1981";
		wait for Clk_period;
		Addr <=  "0011001010011";
		Trees_din <= x"05f3e604";
		wait for Clk_period;
		Addr <=  "0011001010100";
		Trees_din <= x"004b1981";
		wait for Clk_period;
		Addr <=  "0011001010101";
		Trees_din <= x"fff01981";
		wait for Clk_period;
		Addr <=  "0011001010110";
		Trees_din <= x"05f66808";
		wait for Clk_period;
		Addr <=  "0011001010111";
		Trees_din <= x"13039e04";
		wait for Clk_period;
		Addr <=  "0011001011000";
		Trees_din <= x"00b71981";
		wait for Clk_period;
		Addr <=  "0011001011001";
		Trees_din <= x"00291981";
		wait for Clk_period;
		Addr <=  "0011001011010";
		Trees_din <= x"00035a04";
		wait for Clk_period;
		Addr <=  "0011001011011";
		Trees_din <= x"00291981";
		wait for Clk_period;
		Addr <=  "0011001011100";
		Trees_din <= x"ffb61981";
		wait for Clk_period;
		Addr <=  "0011001011101";
		Trees_din <= x"00006604";
		wait for Clk_period;
		Addr <=  "0011001011110";
		Trees_din <= x"001c1981";
		wait for Clk_period;
		Addr <=  "0011001011111";
		Trees_din <= x"007b1981";
		wait for Clk_period;
		Addr <=  "0011001100000";
		Trees_din <= x"1400d108";
		wait for Clk_period;
		Addr <=  "0011001100001";
		Trees_din <= x"020bce04";
		wait for Clk_period;
		Addr <=  "0011001100010";
		Trees_din <= x"ff741a4d";
		wait for Clk_period;
		Addr <=  "0011001100011";
		Trees_din <= x"00251a4d";
		wait for Clk_period;
		Addr <=  "0011001100100";
		Trees_din <= x"020a3130";
		wait for Clk_period;
		Addr <=  "0011001100101";
		Trees_din <= x"1200851c";
		wait for Clk_period;
		Addr <=  "0011001100110";
		Trees_din <= x"1af94c0c";
		wait for Clk_period;
		Addr <=  "0011001100111";
		Trees_din <= x"000b7d08";
		wait for Clk_period;
		Addr <=  "0011001101000";
		Trees_din <= x"07feb504";
		wait for Clk_period;
		Addr <=  "0011001101001";
		Trees_din <= x"00c51a4d";
		wait for Clk_period;
		Addr <=  "0011001101010";
		Trees_din <= x"ffcf1a4d";
		wait for Clk_period;
		Addr <=  "0011001101011";
		Trees_din <= x"ffa31a4d";
		wait for Clk_period;
		Addr <=  "0011001101100";
		Trees_din <= x"0c00b908";
		wait for Clk_period;
		Addr <=  "0011001101101";
		Trees_din <= x"0600b704";
		wait for Clk_period;
		Addr <=  "0011001101110";
		Trees_din <= x"000c1a4d";
		wait for Clk_period;
		Addr <=  "0011001101111";
		Trees_din <= x"ffdf1a4d";
		wait for Clk_period;
		Addr <=  "0011001110000";
		Trees_din <= x"05f54d04";
		wait for Clk_period;
		Addr <=  "0011001110001";
		Trees_din <= x"ff781a4d";
		wait for Clk_period;
		Addr <=  "0011001110010";
		Trees_din <= x"ffe11a4d";
		wait for Clk_period;
		Addr <=  "0011001110011";
		Trees_din <= x"1af94c04";
		wait for Clk_period;
		Addr <=  "0011001110100";
		Trees_din <= x"ff691a4d";
		wait for Clk_period;
		Addr <=  "0011001110101";
		Trees_din <= x"1101b808";
		wait for Clk_period;
		Addr <=  "0011001110110";
		Trees_din <= x"03f95504";
		wait for Clk_period;
		Addr <=  "0011001110111";
		Trees_din <= x"ffd61a4d";
		wait for Clk_period;
		Addr <=  "0011001111000";
		Trees_din <= x"004b1a4d";
		wait for Clk_period;
		Addr <=  "0011001111001";
		Trees_din <= x"0b007f04";
		wait for Clk_period;
		Addr <=  "0011001111010";
		Trees_din <= x"ff8a1a4d";
		wait for Clk_period;
		Addr <=  "0011001111011";
		Trees_din <= x"008e1a4d";
		wait for Clk_period;
		Addr <=  "0011001111100";
		Trees_din <= x"06ff3118";
		wait for Clk_period;
		Addr <=  "0011001111101";
		Trees_din <= x"1c02670c";
		wait for Clk_period;
		Addr <=  "0011001111110";
		Trees_din <= x"020ad304";
		wait for Clk_period;
		Addr <=  "0011001111111";
		Trees_din <= x"ff8d1a4d";
		wait for Clk_period;
		Addr <=  "0011010000000";
		Trees_din <= x"1100d304";
		wait for Clk_period;
		Addr <=  "0011010000001";
		Trees_din <= x"00481a4d";
		wait for Clk_period;
		Addr <=  "0011010000010";
		Trees_din <= x"ffe81a4d";
		wait for Clk_period;
		Addr <=  "0011010000011";
		Trees_din <= x"1403f908";
		wait for Clk_period;
		Addr <=  "0011010000100";
		Trees_din <= x"18016704";
		wait for Clk_period;
		Addr <=  "0011010000101";
		Trees_din <= x"00d41a4d";
		wait for Clk_period;
		Addr <=  "0011010000110";
		Trees_din <= x"003e1a4d";
		wait for Clk_period;
		Addr <=  "0011010000111";
		Trees_din <= x"fffd1a4d";
		wait for Clk_period;
		Addr <=  "0011010001000";
		Trees_din <= x"0e004b10";
		wait for Clk_period;
		Addr <=  "0011010001001";
		Trees_din <= x"0f000208";
		wait for Clk_period;
		Addr <=  "0011010001010";
		Trees_din <= x"01fc5404";
		wait for Clk_period;
		Addr <=  "0011010001011";
		Trees_din <= x"ffce1a4d";
		wait for Clk_period;
		Addr <=  "0011010001100";
		Trees_din <= x"00741a4d";
		wait for Clk_period;
		Addr <=  "0011010001101";
		Trees_din <= x"0b006c04";
		wait for Clk_period;
		Addr <=  "0011010001110";
		Trees_din <= x"00461a4d";
		wait for Clk_period;
		Addr <=  "0011010001111";
		Trees_din <= x"ffe81a4d";
		wait for Clk_period;
		Addr <=  "0011010010000";
		Trees_din <= x"10005304";
		wait for Clk_period;
		Addr <=  "0011010010001";
		Trees_din <= x"ff421a4d";
		wait for Clk_period;
		Addr <=  "0011010010010";
		Trees_din <= x"00271a4d";
		wait for Clk_period;
		Addr <=  "0011010010011";
		Trees_din <= x"0200ea04";
		wait for Clk_period;
		Addr <=  "0011010010100";
		Trees_din <= x"ff8c1aa9";
		wait for Clk_period;
		Addr <=  "0011010010101";
		Trees_din <= x"0b005104";
		wait for Clk_period;
		Addr <=  "0011010010110";
		Trees_din <= x"ff941aa9";
		wait for Clk_period;
		Addr <=  "0011010010111";
		Trees_din <= x"0b005408";
		wait for Clk_period;
		Addr <=  "0011010011000";
		Trees_din <= x"04ff6d04";
		wait for Clk_period;
		Addr <=  "0011010011001";
		Trees_din <= x"00e11aa9";
		wait for Clk_period;
		Addr <=  "0011010011010";
		Trees_din <= x"ffba1aa9";
		wait for Clk_period;
		Addr <=  "0011010011011";
		Trees_din <= x"15004e10";
		wait for Clk_period;
		Addr <=  "0011010011100";
		Trees_din <= x"0c007f08";
		wait for Clk_period;
		Addr <=  "0011010011101";
		Trees_din <= x"1b024804";
		wait for Clk_period;
		Addr <=  "0011010011110";
		Trees_din <= x"ffcd1aa9";
		wait for Clk_period;
		Addr <=  "0011010011111";
		Trees_din <= x"006f1aa9";
		wait for Clk_period;
		Addr <=  "0011010100000";
		Trees_din <= x"0c009604";
		wait for Clk_period;
		Addr <=  "0011010100001";
		Trees_din <= x"ffd81aa9";
		wait for Clk_period;
		Addr <=  "0011010100010";
		Trees_din <= x"000a1aa9";
		wait for Clk_period;
		Addr <=  "0011010100011";
		Trees_din <= x"08003e08";
		wait for Clk_period;
		Addr <=  "0011010100100";
		Trees_din <= x"1600a704";
		wait for Clk_period;
		Addr <=  "0011010100101";
		Trees_din <= x"004f1aa9";
		wait for Clk_period;
		Addr <=  "0011010100110";
		Trees_din <= x"ff9d1aa9";
		wait for Clk_period;
		Addr <=  "0011010100111";
		Trees_din <= x"020b4004";
		wait for Clk_period;
		Addr <=  "0011010101000";
		Trees_din <= x"ff801aa9";
		wait for Clk_period;
		Addr <=  "0011010101001";
		Trees_din <= x"004a1aa9";
		wait for Clk_period;
		Addr <=  "0011010101010";
		Trees_din <= x"0000001f";
		wait for Clk_period;

        -- Reset valid flag
        Valid_node <= '0';
        wait for Clk_period; 
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001010010011010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011100110001";
        wait for Clk_period; 
        Features_din <= "1111100110100001";
        wait for Clk_period; 
        Features_din <= "1111000101100110";
        wait for Clk_period; 
        Features_din <= "0000000111110000";
        wait for Clk_period; 
        Features_din <= "1111010110000110";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "1111110110001001";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000000011001010";
        wait for Clk_period; 
        Features_din <= "0000001000111010";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000011001011";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111100001111000";
        wait for Clk_period; 
        Features_din <= "0000000100110010";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111101100010100";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011011000101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000110011100001";
        wait for Clk_period; 
        Features_din <= "0000000110100110";
        wait for Clk_period; 
        Features_din <= "1111010001011111";
        wait for Clk_period; 
        Features_din <= "1111100100101101";
        wait for Clk_period; 
        Features_din <= "1111011101111111";
        wait for Clk_period; 
        Features_din <= "0000000110110101";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "0000000011000110";
        wait for Clk_period; 
        Features_din <= "0000001001010010";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000100001111";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "0000001100010101";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "1111100000001111";
        wait for Clk_period; 
        Features_din <= "0000000110101100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101110101011";
        wait for Clk_period; 
        Features_din <= "0000001001110101";
        wait for Clk_period; 
        Features_din <= "0000001001110101";
        wait for Clk_period; 
        Features_din <= "0000001001110101";
        wait for Clk_period; 
        Features_din <= "0000001001110101";
        wait for Clk_period; 
        Features_din <= "0000001001110101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000101011110000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000111010001111";
        wait for Clk_period; 
        Features_din <= "0000110000001001";
        wait for Clk_period; 
        Features_din <= "1111011010010100";
        wait for Clk_period; 
        Features_din <= "0000010100100111";
        wait for Clk_period; 
        Features_din <= "1111001001000001";
        wait for Clk_period; 
        Features_din <= "1111101110010001";
        wait for Clk_period; 
        Features_din <= "1111101111110111";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000000011110010";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000100010110";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000011100000";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "1111101000111000";
        wait for Clk_period; 
        Features_din <= "0000000100000110";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "1111100100101010";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(6, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111111011110100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000101010100000";
        wait for Clk_period; 
        Features_din <= "1111100101100111";
        wait for Clk_period; 
        Features_din <= "1111100100101011";
        wait for Clk_period; 
        Features_din <= "1111100000001101";
        wait for Clk_period; 
        Features_din <= "0000010100011000";
        wait for Clk_period; 
        Features_din <= "1111101110010011";
        wait for Clk_period; 
        Features_din <= "1111111100001111";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000010101100";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111011101001110";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110011111110";
        wait for Clk_period; 
        Features_din <= "0000001001010111";
        wait for Clk_period; 
        Features_din <= "0000001001010111";
        wait for Clk_period; 
        Features_din <= "0000001001010111";
        wait for Clk_period; 
        Features_din <= "0000001001010111";
        wait for Clk_period; 
        Features_din <= "0000001001010111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000110101010000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010111011010";
        wait for Clk_period; 
        Features_din <= "0000100011111110";
        wait for Clk_period; 
        Features_din <= "1111011111100001";
        wait for Clk_period; 
        Features_din <= "0000011000000101";
        wait for Clk_period; 
        Features_din <= "1111010101111110";
        wait for Clk_period; 
        Features_din <= "1111110101111101";
        wait for Clk_period; 
        Features_din <= "1111011111110110";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000011111000";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "1111011101110010";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111110010110110";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000110010100011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000100000000001";
        wait for Clk_period; 
        Features_din <= "0000010110000000";
        wait for Clk_period; 
        Features_din <= "1111001101111100";
        wait for Clk_period; 
        Features_din <= "1111101011010101";
        wait for Clk_period; 
        Features_din <= "1111011100000111";
        wait for Clk_period; 
        Features_din <= "0000010100010111";
        wait for Clk_period; 
        Features_din <= "0000000011000010";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000011011111";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000001011111100";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000001010011010";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111100001001010";
        wait for Clk_period; 
        Features_din <= "0000001000101010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101101010011";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000100110000011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000111101010010";
        wait for Clk_period; 
        Features_din <= "0000001011011111";
        wait for Clk_period; 
        Features_din <= "1111101100000110";
        wait for Clk_period; 
        Features_din <= "1111111000111111";
        wait for Clk_period; 
        Features_din <= "1111010001001001";
        wait for Clk_period; 
        Features_din <= "1111110001000111";
        wait for Clk_period; 
        Features_din <= "0000000111100101";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000011011111";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000011000101";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000110000110";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111011110011000";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110001101111";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111110001101000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1110011101100110";
        wait for Clk_period; 
        Features_din <= "0001100010011010";
        wait for Clk_period; 
        Features_din <= "1110011001101100";
        wait for Clk_period; 
        Features_din <= "1111101000101110";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0001001111111111";
        wait for Clk_period; 
        Features_din <= "1111110100000100";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "1111011111101111";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101111011101";
        wait for Clk_period; 
        Features_din <= "0000001001110001";
        wait for Clk_period; 
        Features_din <= "0000001001110001";
        wait for Clk_period; 
        Features_din <= "0000001001110001";
        wait for Clk_period; 
        Features_din <= "0000001001110001";
        wait for Clk_period; 
        Features_din <= "0000001001110001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000010110001011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000101101000011";
        wait for Clk_period; 
        Features_din <= "0000100000110010";
        wait for Clk_period; 
        Features_din <= "1111100111001111";
        wait for Clk_period; 
        Features_din <= "1111101111000110";
        wait for Clk_period; 
        Features_din <= "1111010011101101";
        wait for Clk_period; 
        Features_din <= "1111101101110110";
        wait for Clk_period; 
        Features_din <= "1111101111001110";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000011111011";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "0000000111000100";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000001001001000";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000001011000101";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "1111100001000111";
        wait for Clk_period; 
        Features_din <= "0000000011110001";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111101101011000";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001110110111001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111011000011001";
        wait for Clk_period; 
        Features_din <= "0000110111100111";
        wait for Clk_period; 
        Features_din <= "1111000001100001";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "1111101010100010";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "1111101100101000";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "1111011100110100";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110100110101";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001001101010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000110100100011";
        wait for Clk_period; 
        Features_din <= "0000100011111100";
        wait for Clk_period; 
        Features_din <= "1111101001111010";
        wait for Clk_period; 
        Features_din <= "1111101001000010";
        wait for Clk_period; 
        Features_din <= "1111010101001000";
        wait for Clk_period; 
        Features_din <= "1111110110011101";
        wait for Clk_period; 
        Features_din <= "0000010101000011";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000011011011";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000001011111010";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001010001010";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000110011010";
        wait for Clk_period; 
        Features_din <= "0000000011001110";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "1111111011111110";
        wait for Clk_period; 
        Features_din <= "0000010011011000";
        wait for Clk_period; 
        Features_din <= "1111110110010111";
        wait for Clk_period; 
        Features_din <= "1111110100101010";
        wait for Clk_period; 
        Features_din <= "0000010111011101";
        wait for Clk_period; 
        Features_din <= "1111100111110001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000010010100001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010010111011";
        wait for Clk_period; 
        Features_din <= "0000000110110110";
        wait for Clk_period; 
        Features_din <= "1111100001110101";
        wait for Clk_period; 
        Features_din <= "1111110101110110";
        wait for Clk_period; 
        Features_din <= "1111010110100101";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000010011011101";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000100000000";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111011100000111";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110110011110";
        wait for Clk_period; 
        Features_din <= "0000001001000101";
        wait for Clk_period; 
        Features_din <= "0000001001000101";
        wait for Clk_period; 
        Features_din <= "0000001001000101";
        wait for Clk_period; 
        Features_din <= "0000001001000101";
        wait for Clk_period; 
        Features_din <= "0000001001000101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000010001110111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000100100111111";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111100110100011";
        wait for Clk_period; 
        Features_din <= "1111110100111000";
        wait for Clk_period; 
        Features_din <= "1111100101110100";
        wait for Clk_period; 
        Features_din <= "0000001011001101";
        wait for Clk_period; 
        Features_din <= "1111110110000101";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010110010";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "1111011101011000";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110011101010";
        wait for Clk_period; 
        Features_din <= "0000001001011001";
        wait for Clk_period; 
        Features_din <= "0000001001011001";
        wait for Clk_period; 
        Features_din <= "0000001001011001";
        wait for Clk_period; 
        Features_din <= "0000001001011001";
        wait for Clk_period; 
        Features_din <= "0000001001011001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000110010010111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001000000101110";
        wait for Clk_period; 
        Features_din <= "0000100111100101";
        wait for Clk_period; 
        Features_din <= "1111100000110101";
        wait for Clk_period; 
        Features_din <= "1111111111001011";
        wait for Clk_period; 
        Features_din <= "1111010000110010";
        wait for Clk_period; 
        Features_din <= "0000010101001111";
        wait for Clk_period; 
        Features_din <= "1111010010111000";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000011101100";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000100000111";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "1111011110010010";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111110001111100";
        wait for Clk_period; 
        Features_din <= "0000001001100100";
        wait for Clk_period; 
        Features_din <= "0000001001100100";
        wait for Clk_period; 
        Features_din <= "0000001001100100";
        wait for Clk_period; 
        Features_din <= "0000001001100100";
        wait for Clk_period; 
        Features_din <= "0000001001100100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000010110011010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111001011100001";
        wait for Clk_period; 
        Features_din <= "0001010010100000";
        wait for Clk_period; 
        Features_din <= "1111001011011111";
        wait for Clk_period; 
        Features_din <= "0000110100000110";
        wait for Clk_period; 
        Features_din <= "1111101101110110";
        wait for Clk_period; 
        Features_din <= "1111101000100100";
        wait for Clk_period; 
        Features_din <= "1111011010101101";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000011011111";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000011101010";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "1111011011101100";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110111100001";
        wait for Clk_period; 
        Features_din <= "0000001000111101";
        wait for Clk_period; 
        Features_din <= "0000001000111101";
        wait for Clk_period; 
        Features_din <= "0000001000111101";
        wait for Clk_period; 
        Features_din <= "0000001000111101";
        wait for Clk_period; 
        Features_din <= "0000001000111101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001000001001001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001001100110110";
        wait for Clk_period; 
        Features_din <= "0000000011000111";
        wait for Clk_period; 
        Features_din <= "1111001000001010";
        wait for Clk_period; 
        Features_din <= "1111110000101010";
        wait for Clk_period; 
        Features_din <= "1111000011110101";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "1111010111010110";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "0000001000101010";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "0000001001010010";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111011101000010";
        wait for Clk_period; 
        Features_din <= "0000000011111010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110100011001";
        wait for Clk_period; 
        Features_din <= "0000001001010100";
        wait for Clk_period; 
        Features_din <= "0000001001010100";
        wait for Clk_period; 
        Features_din <= "0000001001010100";
        wait for Clk_period; 
        Features_din <= "0000001001010100";
        wait for Clk_period; 
        Features_din <= "0000001001010100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000010000101110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000110000110010";
        wait for Clk_period; 
        Features_din <= "0000010101111011";
        wait for Clk_period; 
        Features_din <= "1111010111001101";
        wait for Clk_period; 
        Features_din <= "1111111000010010";
        wait for Clk_period; 
        Features_din <= "1111011000000001";
        wait for Clk_period; 
        Features_din <= "1111111110100000";
        wait for Clk_period; 
        Features_din <= "1111110101101100";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000011100010";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "0000000100001011";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000011110011";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111011111010111";
        wait for Clk_period; 
        Features_din <= "0000000011001100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110000000011";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111100011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000100110100110";
        wait for Clk_period; 
        Features_din <= "0000011010001101";
        wait for Clk_period; 
        Features_din <= "1111101001011101";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "1111101000001101";
        wait for Clk_period; 
        Features_din <= "1111111001011101";
        wait for Clk_period; 
        Features_din <= "1111111011001101";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000011101100";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000110011110";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "1111100000101110";
        wait for Clk_period; 
        Features_din <= "0000000011100111";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111101101111011";
        wait for Clk_period; 
        Features_din <= "0000001001111000";
        wait for Clk_period; 
        Features_din <= "0000001001111000";
        wait for Clk_period; 
        Features_din <= "0000001001111000";
        wait for Clk_period; 
        Features_din <= "0000001001111000";
        wait for Clk_period; 
        Features_din <= "0000001001111000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001100101001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111011110101010";
        wait for Clk_period; 
        Features_din <= "0000011100001001";
        wait for Clk_period; 
        Features_din <= "1111001011011000";
        wait for Clk_period; 
        Features_din <= "1111111111110000";
        wait for Clk_period; 
        Features_din <= "1111100011111100";
        wait for Clk_period; 
        Features_din <= "0001110000000001";
        wait for Clk_period; 
        Features_din <= "1111011100011000";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000100000011";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "1111011110000010";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110010011000";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000101110100010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000110101101001";
        wait for Clk_period; 
        Features_din <= "0000011011111101";
        wait for Clk_period; 
        Features_din <= "1111101010001100";
        wait for Clk_period; 
        Features_din <= "0000011110110001";
        wait for Clk_period; 
        Features_din <= "1111001101010001";
        wait for Clk_period; 
        Features_din <= "1111111000110001";
        wait for Clk_period; 
        Features_din <= "1111011101001101";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000011100101";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000011101110";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "1111011110011000";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110001101111";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001101001011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000101100101010";
        wait for Clk_period; 
        Features_din <= "0000100000010100";
        wait for Clk_period; 
        Features_din <= "1111010100010011";
        wait for Clk_period; 
        Features_din <= "0000001000111110";
        wait for Clk_period; 
        Features_din <= "1111010101100101";
        wait for Clk_period; 
        Features_din <= "0000010010110001";
        wait for Clk_period; 
        Features_din <= "1111110010010111";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000011110010";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "1111011101001110";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111110011111111";
        wait for Clk_period; 
        Features_din <= "0000001001010111";
        wait for Clk_period; 
        Features_din <= "0000001001010111";
        wait for Clk_period; 
        Features_din <= "0000001001010111";
        wait for Clk_period; 
        Features_din <= "0000001001010111";
        wait for Clk_period; 
        Features_din <= "0000001001010111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001000110100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000110001111101";
        wait for Clk_period; 
        Features_din <= "1111011000011100";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "0000000011011110";
        wait for Clk_period; 
        Features_din <= "1111011010101011";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "0000000110100000";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000001001010011";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000001011010010";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111011100111110";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110100100010";
        wait for Clk_period; 
        Features_din <= "0000001001010011";
        wait for Clk_period; 
        Features_din <= "0000001001010011";
        wait for Clk_period; 
        Features_din <= "0000001001010011";
        wait for Clk_period; 
        Features_din <= "0000001001010011";
        wait for Clk_period; 
        Features_din <= "0000001001010011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000111011110111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000110010110110";
        wait for Clk_period; 
        Features_din <= "0000011100110101";
        wait for Clk_period; 
        Features_din <= "1111010111111111";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "1111000101011110";
        wait for Clk_period; 
        Features_din <= "0000010010010010";
        wait for Clk_period; 
        Features_din <= "1111010011001011";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000011100001";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000011001110";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000101101110";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111100001101011";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111101100100101";
        wait for Clk_period; 
        Features_din <= "0000001001111101";
        wait for Clk_period; 
        Features_din <= "0000001001111101";
        wait for Clk_period; 
        Features_din <= "0000001001111101";
        wait for Clk_period; 
        Features_din <= "0000001001111101";
        wait for Clk_period; 
        Features_din <= "0000001001111101";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000100101000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100001011";
        wait for Clk_period; 
        Features_din <= "0000100000100000";
        wait for Clk_period; 
        Features_din <= "0001010101001001";
        wait for Clk_period; 
        Features_din <= "1111010010001000";
        wait for Clk_period; 
        Features_din <= "1111101100001011";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111110111001001";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000011100111";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000011000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000101010111";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111011110100001";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110001100000";
        wait for Clk_period; 
        Features_din <= "0000001001100110";
        wait for Clk_period; 
        Features_din <= "0000001001100110";
        wait for Clk_period; 
        Features_din <= "0000001001100110";
        wait for Clk_period; 
        Features_din <= "0000001001100110";
        wait for Clk_period; 
        Features_din <= "0000001001100110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(6, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111110010101111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000100010000011";
        wait for Clk_period; 
        Features_din <= "0000011010010010";
        wait for Clk_period; 
        Features_din <= "1111101101011001";
        wait for Clk_period; 
        Features_din <= "1111101111010100";
        wait for Clk_period; 
        Features_din <= "0000000011010110";
        wait for Clk_period; 
        Features_din <= "1111110000101001";
        wait for Clk_period; 
        Features_din <= "0000001100101001";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000011111100";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000011100011";
        wait for Clk_period; 
        Features_din <= "0000000011101100";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "1111100001001000";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101101010110";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000100010111110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010111100111";
        wait for Clk_period; 
        Features_din <= "0000010111001101";
        wait for Clk_period; 
        Features_din <= "1111001100110100";
        wait for Clk_period; 
        Features_din <= "1111101100000110";
        wait for Clk_period; 
        Features_din <= "1111100000111010";
        wait for Clk_period; 
        Features_din <= "0000100110100101";
        wait for Clk_period; 
        Features_din <= "1111101110100100";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000011100001";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000101101001";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111100011000000";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111101010110101";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011001000001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001001011111";
        wait for Clk_period; 
        Features_din <= "0000001010101111";
        wait for Clk_period; 
        Features_din <= "1111100011001010";
        wait for Clk_period; 
        Features_din <= "1111100110100100";
        wait for Clk_period; 
        Features_din <= "0000101001101100";
        wait for Clk_period; 
        Features_din <= "0000011010001001";
        wait for Clk_period; 
        Features_din <= "1111110010111000";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000011100100";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "1111011111001101";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111110000010101";
        wait for Clk_period; 
        Features_din <= "0000001001101101";
        wait for Clk_period; 
        Features_din <= "0000001001101101";
        wait for Clk_period; 
        Features_din <= "0000001001101101";
        wait for Clk_period; 
        Features_din <= "0000001001101101";
        wait for Clk_period; 
        Features_din <= "0000001001101101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011101100001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000111001001000";
        wait for Clk_period; 
        Features_din <= "0000010110011100";
        wait for Clk_period; 
        Features_din <= "1111101000101011";
        wait for Clk_period; 
        Features_din <= "0000001011011010";
        wait for Clk_period; 
        Features_din <= "1111011110011011";
        wait for Clk_period; 
        Features_din <= "1111101110011011";
        wait for Clk_period; 
        Features_din <= "1111100100100111";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000011011110";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000000011000110";
        wait for Clk_period; 
        Features_din <= "0000000011101010";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000011011101";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "1111011110001000";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110010001110";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011001011111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001000010001010";
        wait for Clk_period; 
        Features_din <= "0000100100010110";
        wait for Clk_period; 
        Features_din <= "1111000001011110";
        wait for Clk_period; 
        Features_din <= "1111101011001100";
        wait for Clk_period; 
        Features_din <= "1111000000000010";
        wait for Clk_period; 
        Features_din <= "0001000100110110";
        wait for Clk_period; 
        Features_din <= "1111100011111111";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000000011001000";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000110111110";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "1111100010111110";
        wait for Clk_period; 
        Features_din <= "0000000101011111";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111101010111001";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001001011111100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000110010010111";
        wait for Clk_period; 
        Features_din <= "0000101110100000";
        wait for Clk_period; 
        Features_din <= "1111011101101111";
        wait for Clk_period; 
        Features_din <= "0000010100000111";
        wait for Clk_period; 
        Features_din <= "1111010110000111";
        wait for Clk_period; 
        Features_din <= "0000000011000101";
        wait for Clk_period; 
        Features_din <= "1111010011111010";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000011101000";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000100111001";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "1111011110111001";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111110000110110";
        wait for Clk_period; 
        Features_din <= "0000001001101010";
        wait for Clk_period; 
        Features_din <= "0000001001101010";
        wait for Clk_period; 
        Features_din <= "0000001001101010";
        wait for Clk_period; 
        Features_din <= "0000001001101010";
        wait for Clk_period; 
        Features_din <= "0000001001101010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000111001110011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000101101101100";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "1111001110101001";
        wait for Clk_period; 
        Features_din <= "0000000110100111";
        wait for Clk_period; 
        Features_din <= "1111001110111001";
        wait for Clk_period; 
        Features_din <= "1111111000000000";
        wait for Clk_period; 
        Features_din <= "1111101101110001";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "1111011110101100";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111110001001100";
        wait for Clk_period; 
        Features_din <= "0000001001101000";
        wait for Clk_period; 
        Features_din <= "0000001001101000";
        wait for Clk_period; 
        Features_din <= "0000001001101000";
        wait for Clk_period; 
        Features_din <= "0000001001101000";
        wait for Clk_period; 
        Features_din <= "0000001001101000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010101001111100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100011100";
        wait for Clk_period; 
        Features_din <= "0000110100001100";
        wait for Clk_period; 
        Features_din <= "1110111001101111";
        wait for Clk_period; 
        Features_din <= "0001010010011111";
        wait for Clk_period; 
        Features_din <= "1111010111011001";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "1110111101100111";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000100011101";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000101110101";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111100000110011";
        wait for Clk_period; 
        Features_din <= "0000000010111101";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111101101110100";
        wait for Clk_period; 
        Features_din <= "0000001001111000";
        wait for Clk_period; 
        Features_din <= "0000001001111000";
        wait for Clk_period; 
        Features_din <= "0000001001111000";
        wait for Clk_period; 
        Features_din <= "0000001001111000";
        wait for Clk_period; 
        Features_din <= "0000001001111000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000100010110000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000111011111011";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "1111110001001111";
        wait for Clk_period; 
        Features_din <= "1111100101010010";
        wait for Clk_period; 
        Features_din <= "1111011010110011";
        wait for Clk_period; 
        Features_din <= "1111101111000101";
        wait for Clk_period; 
        Features_din <= "1111101101010100";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "0000001010100110";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000001000000110";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000001000110111";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "1111011101011111";
        wait for Clk_period; 
        Features_din <= "0000000101000101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110011011100";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000010101001010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1110111010100010";
        wait for Clk_period; 
        Features_din <= "0000100011010010";
        wait for Clk_period; 
        Features_din <= "1111011011001010";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "0000000110001010";
        wait for Clk_period; 
        Features_din <= "0001001010000000";
        wait for Clk_period; 
        Features_din <= "1111110010110100";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000011110000";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "1111011110010011";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110001111010";
        wait for Clk_period; 
        Features_din <= "0000001001100100";
        wait for Clk_period; 
        Features_din <= "0000001001100100";
        wait for Clk_period; 
        Features_din <= "0000001001100100";
        wait for Clk_period; 
        Features_din <= "0000001001100100";
        wait for Clk_period; 
        Features_din <= "0000001001100100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001011001101011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000011110001111";
        wait for Clk_period; 
        Features_din <= "1111100110100011";
        wait for Clk_period; 
        Features_din <= "0000100011011001";
        wait for Clk_period; 
        Features_din <= "1111110000101000";
        wait for Clk_period; 
        Features_din <= "1111111111011100";
        wait for Clk_period; 
        Features_din <= "1111101100100011";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000011011011";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000011000010";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000100010011";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111100001001000";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111101101010110";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(3, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111101100100001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011000010011";
        wait for Clk_period; 
        Features_din <= "0000101110110001";
        wait for Clk_period; 
        Features_din <= "0001001110110001";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111100111110011";
        wait for Clk_period; 
        Features_din <= "1111100110011101";
        wait for Clk_period; 
        Features_din <= "1111101111100110";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "0000000101010010";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000010111";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "1111011101011110";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110011011110";
        wait for Clk_period; 
        Features_din <= "0000001001011010";
        wait for Clk_period; 
        Features_din <= "0000001001011010";
        wait for Clk_period; 
        Features_din <= "0000001001011010";
        wait for Clk_period; 
        Features_din <= "0000001001011010";
        wait for Clk_period; 
        Features_din <= "0000001001011010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(6, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111110010001100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001000001101";
        wait for Clk_period; 
        Features_din <= "1111101111010000";
        wait for Clk_period; 
        Features_din <= "1111010000010001";
        wait for Clk_period; 
        Features_din <= "1111010110101001";
        wait for Clk_period; 
        Features_din <= "0001000001110000";
        wait for Clk_period; 
        Features_din <= "0000100100101111";
        wait for Clk_period; 
        Features_din <= "0000001011010110";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000000011001000";
        wait for Clk_period; 
        Features_din <= "0000000101000001";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000110100011";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "1111100011000011";
        wait for Clk_period; 
        Features_din <= "0000000100010111";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "1111101010110011";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000100111110011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111100001101010";
        wait for Clk_period; 
        Features_din <= "0000111101001011";
        wait for Clk_period; 
        Features_din <= "1111111011110011";
        wait for Clk_period; 
        Features_din <= "1111111110100010";
        wait for Clk_period; 
        Features_din <= "0000101011110011";
        wait for Clk_period; 
        Features_din <= "0000001011010000";
        wait for Clk_period; 
        Features_din <= "1111101000011000";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000011010010";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000011100101";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000101001101";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "1111011111000110";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110000100000";
        wait for Clk_period; 
        Features_din <= "0000001001101100";
        wait for Clk_period; 
        Features_din <= "0000001001101100";
        wait for Clk_period; 
        Features_din <= "0000001001101100";
        wait for Clk_period; 
        Features_din <= "0000001001101100";
        wait for Clk_period; 
        Features_din <= "0000001001101100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011000010111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000100101001111";
        wait for Clk_period; 
        Features_din <= "0000011001110000";
        wait for Clk_period; 
        Features_din <= "1111011000100000";
        wait for Clk_period; 
        Features_din <= "1111110101000111";
        wait for Clk_period; 
        Features_din <= "1111100010001010";
        wait for Clk_period; 
        Features_din <= "1111110011010010";
        wait for Clk_period; 
        Features_din <= "1111111101011100";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000011110111";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000000100011001";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000111000110";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001100010111";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000110001110";
        wait for Clk_period; 
        Features_din <= "0000001000111110";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "1111111010001011";
        wait for Clk_period; 
        Features_din <= "0000010010110110";
        wait for Clk_period; 
        Features_din <= "1111110101100110";
        wait for Clk_period; 
        Features_din <= "1111110101100010";
        wait for Clk_period; 
        Features_din <= "0000011000110000";
        wait for Clk_period; 
        Features_din <= "1111101000111010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011100111000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000110000001000";
        wait for Clk_period; 
        Features_din <= "1111011010010111";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "1111001011010001";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "1111110011111001";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000011111000";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000010010001";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000100001110";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "1111011101110110";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110010101111";
        wait for Clk_period; 
        Features_din <= "0000001001011111";
        wait for Clk_period; 
        Features_din <= "0000001001011111";
        wait for Clk_period; 
        Features_din <= "0000001001011111";
        wait for Clk_period; 
        Features_din <= "0000001001011111";
        wait for Clk_period; 
        Features_din <= "0000001001011111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000010110101001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000110100111110";
        wait for Clk_period; 
        Features_din <= "0000001011101110";
        wait for Clk_period; 
        Features_din <= "1111100100101111";
        wait for Clk_period; 
        Features_din <= "1111101001001101";
        wait for Clk_period; 
        Features_din <= "1111010010000011";
        wait for Clk_period; 
        Features_din <= "1111110001000000";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111011101110001";
        wait for Clk_period; 
        Features_din <= "0000000000101000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110010111001";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000010001110001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011110010011";
        wait for Clk_period; 
        Features_din <= "0000101011010111";
        wait for Clk_period; 
        Features_din <= "1111111000010000";
        wait for Clk_period; 
        Features_din <= "1111111111010001";
        wait for Clk_period; 
        Features_din <= "1111011001011010";
        wait for Clk_period; 
        Features_din <= "0000001011111111";
        wait for Clk_period; 
        Features_din <= "1111110001000001";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000011101010";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000100111001";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111111010010001";
        wait for Clk_period; 
        Features_din <= "0000000100000000";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000001100000010";
        wait for Clk_period; 
        Features_din <= "1111101111010010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000000101111000";
        wait for Clk_period; 
        Features_din <= "1111100100001111";
        wait for Clk_period; 
        Features_din <= "0000010001111101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011001101110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000100101001010";
        wait for Clk_period; 
        Features_din <= "0000100000010011";
        wait for Clk_period; 
        Features_din <= "1111011011110110";
        wait for Clk_period; 
        Features_din <= "1111111010111100";
        wait for Clk_period; 
        Features_din <= "1111011101000000";
        wait for Clk_period; 
        Features_din <= "1111111111110111";
        wait for Clk_period; 
        Features_din <= "1111111101000000";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000011100001";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000011000101";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "0000000000001100";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000100110000";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "1111011110110110";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110000111010";
        wait for Clk_period; 
        Features_din <= "0000001001101001";
        wait for Clk_period; 
        Features_din <= "0000001001101001";
        wait for Clk_period; 
        Features_din <= "0000001001101001";
        wait for Clk_period; 
        Features_din <= "0000001001101001";
        wait for Clk_period; 
        Features_din <= "0000001001101001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000100100100101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111011111011";
        wait for Clk_period; 
        Features_din <= "1111111111111100";
        wait for Clk_period; 
        Features_din <= "1111010000010000";
        wait for Clk_period; 
        Features_din <= "1111101110000101";
        wait for Clk_period; 
        Features_din <= "0000100100100101";
        wait for Clk_period; 
        Features_din <= "0000000011001011";
        wait for Clk_period; 
        Features_din <= "0000010100110100";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000011010000";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000000011101110";
        wait for Clk_period; 
        Features_din <= "0000000101001001";
        wait for Clk_period; 
        Features_din <= "0000000000011111";
        wait for Clk_period; 
        Features_din <= "0000000100101011";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000011110100";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "1111100101110110";
        wait for Clk_period; 
        Features_din <= "0000000101110000";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "1111100111100101";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000100000100101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "0000101000011111";
        wait for Clk_period; 
        Features_din <= "1111011001001001";
        wait for Clk_period; 
        Features_din <= "0000010010001000";
        wait for Clk_period; 
        Features_din <= "1111011010001100";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "1111111111110011";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000011101101";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000011010011";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "1111011101001010";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111110100000111";
        wait for Clk_period; 
        Features_din <= "0000001001010110";
        wait for Clk_period; 
        Features_din <= "0000001001010110";
        wait for Clk_period; 
        Features_din <= "0000001001010110";
        wait for Clk_period; 
        Features_din <= "0000001001010110";
        wait for Clk_period; 
        Features_din <= "0000001001010110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001000000100001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001001101110000";
        wait for Clk_period; 
        Features_din <= "0000101000001000";
        wait for Clk_period; 
        Features_din <= "1111011110010111";
        wait for Clk_period; 
        Features_din <= "0000011101111000";
        wait for Clk_period; 
        Features_din <= "1110110010111110";
        wait for Clk_period; 
        Features_din <= "0000010100011001";
        wait for Clk_period; 
        Features_din <= "1111100111101001";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000001010101101";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000001011110000";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "1111100100100100";
        wait for Clk_period; 
        Features_din <= "0000000100100101";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "1111101000111110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011110010111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000101011101010";
        wait for Clk_period; 
        Features_din <= "0000110011000010";
        wait for Clk_period; 
        Features_din <= "1111101100100010";
        wait for Clk_period; 
        Features_din <= "1111110010100000";
        wait for Clk_period; 
        Features_din <= "1110111111110110";
        wait for Clk_period; 
        Features_din <= "1111101101010010";
        wait for Clk_period; 
        Features_din <= "1111110101000101";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000011011111";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000111111010";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "1111100011010001";
        wait for Clk_period; 
        Features_din <= "0000000100011101";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111101010100001";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000110101010001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111011010111010";
        wait for Clk_period; 
        Features_din <= "0001000100011011";
        wait for Clk_period; 
        Features_din <= "1110100111010100";
        wait for Clk_period; 
        Features_din <= "0000010100110110";
        wait for Clk_period; 
        Features_din <= "1111110000110110";
        wait for Clk_period; 
        Features_din <= "0000100001000111";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000011101001";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000001011011100";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000001011001001";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111100000010101";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111101110100001";
        wait for Clk_period; 
        Features_din <= "0000001001110101";
        wait for Clk_period; 
        Features_din <= "0000001001110101";
        wait for Clk_period; 
        Features_din <= "0000001001110101";
        wait for Clk_period; 
        Features_din <= "0000001001110101";
        wait for Clk_period; 
        Features_din <= "0000001001110101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000111110100010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000111001111111";
        wait for Clk_period; 
        Features_din <= "0000010100111000";
        wait for Clk_period; 
        Features_din <= "1111010000110101";
        wait for Clk_period; 
        Features_din <= "0000010011111011";
        wait for Clk_period; 
        Features_din <= "1111101000010000";
        wait for Clk_period; 
        Features_din <= "0000001000100011";
        wait for Clk_period; 
        Features_din <= "1111011101111111";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000001100001100";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000001010010100";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111100100101110";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111101000110011";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000100100011110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001000101101";
        wait for Clk_period; 
        Features_din <= "0000010100001011";
        wait for Clk_period; 
        Features_din <= "1111001101111000";
        wait for Clk_period; 
        Features_din <= "1111110111111000";
        wait for Clk_period; 
        Features_din <= "1111101001110000";
        wait for Clk_period; 
        Features_din <= "1111101101011111";
        wait for Clk_period; 
        Features_din <= "0000011011000001";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "0000000011010000";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "0000000100000001";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000111010001";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "1111101000101101";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "1111100100110100";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001000110110100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001000110101100";
        wait for Clk_period; 
        Features_din <= "0000100000111001";
        wait for Clk_period; 
        Features_din <= "1111011010101100";
        wait for Clk_period; 
        Features_din <= "1111111100011110";
        wait for Clk_period; 
        Features_din <= "1111001000111111";
        wait for Clk_period; 
        Features_din <= "0000001010001100";
        wait for Clk_period; 
        Features_din <= "1111001000110111";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000011011101";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "0000001000000010";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000101010100";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000001001001111";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000001010010011";
        wait for Clk_period; 
        Features_din <= "0000001100010000";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "1111100101101100";
        wait for Clk_period; 
        Features_din <= "0000001000110100";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "1111100111110000";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001011111100010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111100001101100";
        wait for Clk_period; 
        Features_din <= "0000111100000101";
        wait for Clk_period; 
        Features_din <= "1111010011011000";
        wait for Clk_period; 
        Features_din <= "1111101010111010";
        wait for Clk_period; 
        Features_din <= "1111010110010001";
        wait for Clk_period; 
        Features_din <= "1111110111100000";
        wait for Clk_period; 
        Features_din <= "1111111001001110";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000011011010";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000000011001010";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000101100111";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "1111100001111110";
        wait for Clk_period; 
        Features_din <= "0000000111101100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101100001100";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011000111110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011101011001";
        wait for Clk_period; 
        Features_din <= "0000010011100000";
        wait for Clk_period; 
        Features_din <= "1111100110000101";
        wait for Clk_period; 
        Features_din <= "1111100100100011";
        wait for Clk_period; 
        Features_din <= "1111110011101100";
        wait for Clk_period; 
        Features_din <= "0000011100000011";
        wait for Clk_period; 
        Features_din <= "1111111100010001";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "0000000011011100";
        wait for Clk_period; 
        Features_din <= "0000001001010100";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000001001100110";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000101000111";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000001011111110";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111111011010001";
        wait for Clk_period; 
        Features_din <= "0000001010001101";
        wait for Clk_period; 
        Features_din <= "0000000111100001";
        wait for Clk_period; 
        Features_din <= "1111111111111101";
        wait for Clk_period; 
        Features_din <= "0000001011000101";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "0000000111000111";
        wait for Clk_period; 
        Features_din <= "1111011101010101";
        wait for Clk_period; 
        Features_din <= "0000010011110011";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0010000101010000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111101000110110";
        wait for Clk_period; 
        Features_din <= "0000101110001010";
        wait for Clk_period; 
        Features_din <= "1111010110001001";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "1111010011001101";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "1111100111001000";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000011011101";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000011110001";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000110111111";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000001100001011";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "1111101011001100";
        wait for Clk_period; 
        Features_din <= "0000000101100100";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "1111100010101110";
        wait for Clk_period; 
        Features_din <= "0000001010000001";
        wait for Clk_period; 
        Features_din <= "0000001010000001";
        wait for Clk_period; 
        Features_din <= "0000001010000001";
        wait for Clk_period; 
        Features_din <= "0000001010000001";
        wait for Clk_period; 
        Features_din <= "0000001010000001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000101011110001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011000111001";
        wait for Clk_period; 
        Features_din <= "0000011110001110";
        wait for Clk_period; 
        Features_din <= "1111101101000101";
        wait for Clk_period; 
        Features_din <= "0000110001100000";
        wait for Clk_period; 
        Features_din <= "1111001101111111";
        wait for Clk_period; 
        Features_din <= "0000011010000110";
        wait for Clk_period; 
        Features_din <= "1111110111100101";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "0000001000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000001001100110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "1111100011011100";
        wait for Clk_period; 
        Features_din <= "0000000100101110";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "1111101010010011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000010110010001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001000110100010";
        wait for Clk_period; 
        Features_din <= "0000000110101010";
        wait for Clk_period; 
        Features_din <= "1111100100110101";
        wait for Clk_period; 
        Features_din <= "0000001011000000";
        wait for Clk_period; 
        Features_din <= "1111011001101001";
        wait for Clk_period; 
        Features_din <= "0000010111001100";
        wait for Clk_period; 
        Features_din <= "1111010111100000";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000011101110";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000101101000";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "1111011110000101";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110010010100";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011011101000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000110101101110";
        wait for Clk_period; 
        Features_din <= "0000011001111100";
        wait for Clk_period; 
        Features_din <= "1111101010000001";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "1111010100001101";
        wait for Clk_period; 
        Features_din <= "1111110010001000";
        wait for Clk_period; 
        Features_din <= "1111110100101101";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "1111011111101001";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101111100110";
        wait for Clk_period; 
        Features_din <= "0000001001110000";
        wait for Clk_period; 
        Features_din <= "0000001001110000";
        wait for Clk_period; 
        Features_din <= "0000001001110000";
        wait for Clk_period; 
        Features_din <= "0000001001110000";
        wait for Clk_period; 
        Features_din <= "0000001001110000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111110010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010110000001";
        wait for Clk_period; 
        Features_din <= "0000001000101101";
        wait for Clk_period; 
        Features_din <= "1111100110000100";
        wait for Clk_period; 
        Features_din <= "1111111000011101";
        wait for Clk_period; 
        Features_din <= "1111110001100110";
        wait for Clk_period; 
        Features_din <= "1111110111000101";
        wait for Clk_period; 
        Features_din <= "0000011100010001";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "1111100010000110";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111101100000001";
        wait for Clk_period; 
        Features_din <= "0000001001111111";
        wait for Clk_period; 
        Features_din <= "0000001001111111";
        wait for Clk_period; 
        Features_din <= "0000001001111111";
        wait for Clk_period; 
        Features_din <= "0000001001111111";
        wait for Clk_period; 
        Features_din <= "0000001001111111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000010001011111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000000111011111";
        wait for Clk_period; 
        Features_din <= "0001001100111000";
        wait for Clk_period; 
        Features_din <= "1111101101110101";
        wait for Clk_period; 
        Features_din <= "0000010101001100";
        wait for Clk_period; 
        Features_din <= "1111010001001000";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "1111010100010010";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "0000000111101100";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000011111011";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000000101000001";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "1111101001001111";
        wait for Clk_period; 
        Features_din <= "0000001001001010";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111100100010110";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000101001001110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000110100111100";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "1111011010110101";
        wait for Clk_period; 
        Features_din <= "0000001011000010";
        wait for Clk_period; 
        Features_din <= "1111010010001100";
        wait for Clk_period; 
        Features_din <= "1111111110111011";
        wait for Clk_period; 
        Features_din <= "1111011110111101";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000011100111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000111100011";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111100000011100";
        wait for Clk_period; 
        Features_din <= "0000000010111010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101110010110";
        wait for Clk_period; 
        Features_din <= "0000001001110110";
        wait for Clk_period; 
        Features_din <= "0000001001110110";
        wait for Clk_period; 
        Features_din <= "0000001001110110";
        wait for Clk_period; 
        Features_din <= "0000001001110110";
        wait for Clk_period; 
        Features_din <= "0000001001110110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000110001110110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000111101010001";
        wait for Clk_period; 
        Features_din <= "0000110110110110";
        wait for Clk_period; 
        Features_din <= "1111010101101000";
        wait for Clk_period; 
        Features_din <= "0000001011111100";
        wait for Clk_period; 
        Features_din <= "1110110111010000";
        wait for Clk_period; 
        Features_din <= "1111111111101001";
        wait for Clk_period; 
        Features_din <= "1111011100101110";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000011101110";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000100001011";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "1111011110100010";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110001011110";
        wait for Clk_period; 
        Features_din <= "0000001001100110";
        wait for Clk_period; 
        Features_din <= "0000001001100110";
        wait for Clk_period; 
        Features_din <= "0000001001100110";
        wait for Clk_period; 
        Features_din <= "0000001001100110";
        wait for Clk_period; 
        Features_din <= "0000001001100110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000111000110111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001001011111101";
        wait for Clk_period; 
        Features_din <= "0000011110111100";
        wait for Clk_period; 
        Features_din <= "1111010001011010";
        wait for Clk_period; 
        Features_din <= "1111111011011111";
        wait for Clk_period; 
        Features_din <= "1111001010110111";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111010011101010";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000010101011";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000010111110";
        wait for Clk_period; 
        Features_din <= "0000000111111111";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000001100101101";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "0000000101100010";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "1111011111100110";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101111101011";
        wait for Clk_period; 
        Features_din <= "0000001001110000";
        wait for Clk_period; 
        Features_din <= "0000001001110000";
        wait for Clk_period; 
        Features_din <= "0000001001110000";
        wait for Clk_period; 
        Features_din <= "0000001001110000";
        wait for Clk_period; 
        Features_din <= "0000001001110000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000111011100110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000010110011011";
        wait for Clk_period; 
        Features_din <= "1110110101111101";
        wait for Clk_period; 
        Features_din <= "0000110100011010";
        wait for Clk_period; 
        Features_din <= "1111101010011000";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "1111001000101011";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000010110010";
        wait for Clk_period; 
        Features_din <= "0000001001000111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000100110011";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000001011110111";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000101101011";
        wait for Clk_period; 
        Features_din <= "0000001011110010";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "1111101000001100";
        wait for Clk_period; 
        Features_din <= "0000001001101101";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "1111100101010010";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001000010101101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000101100011010";
        wait for Clk_period; 
        Features_din <= "0000011101000000";
        wait for Clk_period; 
        Features_din <= "1111010011001011";
        wait for Clk_period; 
        Features_din <= "0000001010001011";
        wait for Clk_period; 
        Features_din <= "1111010110110010";
        wait for Clk_period; 
        Features_din <= "0000000101001001";
        wait for Clk_period; 
        Features_din <= "1111001111010011";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000010111000";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000001000001101";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "1111011111100001";
        wait for Clk_period; 
        Features_din <= "0000000011011010";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111101111110010";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001000100010111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000100010100001";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "1111001010110000";
        wait for Clk_period; 
        Features_din <= "1111110100001100";
        wait for Clk_period; 
        Features_din <= "1111110000001110";
        wait for Clk_period; 
        Features_din <= "0000000100111010";
        wait for Clk_period; 
        Features_din <= "1111011010111010";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000011110110";
        wait for Clk_period; 
        Features_din <= "0000001001001100";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000110011011";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "0000001011011011";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111100010111011";
        wait for Clk_period; 
        Features_din <= "0000000111100100";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "1111101010111100";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000001010000010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011101110111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001100100111";
        wait for Clk_period; 
        Features_din <= "0000100111010101";
        wait for Clk_period; 
        Features_din <= "1111100010110110";
        wait for Clk_period; 
        Features_din <= "1111110001101001";
        wait for Clk_period; 
        Features_din <= "1111101110111000";
        wait for Clk_period; 
        Features_din <= "0000010011011000";
        wait for Clk_period; 
        Features_din <= "0000011001101010";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000100000000";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "1111011010111101";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111111001100011";
        wait for Clk_period; 
        Features_din <= "0000001000101101";
        wait for Clk_period; 
        Features_din <= "0000001000101101";
        wait for Clk_period; 
        Features_din <= "0000001000101101";
        wait for Clk_period; 
        Features_din <= "0000001000101101";
        wait for Clk_period; 
        Features_din <= "0000001000101101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001001010110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111010110001";
        wait for Clk_period; 
        Features_din <= "0000110101111001";
        wait for Clk_period; 
        Features_din <= "1111100000000010";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "1111100010001100";
        wait for Clk_period; 
        Features_din <= "0000100001100001";
        wait for Clk_period; 
        Features_din <= "1111110011111011";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000011111001";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "1111011110110011";
        wait for Clk_period; 
        Features_din <= "0000000000011000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110001000001";
        wait for Clk_period; 
        Features_din <= "0000001001101001";
        wait for Clk_period; 
        Features_din <= "0000001001101001";
        wait for Clk_period; 
        Features_din <= "0000001001101001";
        wait for Clk_period; 
        Features_din <= "0000001001101001";
        wait for Clk_period; 
        Features_din <= "0000001001101001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011001111001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000101111110011";
        wait for Clk_period; 
        Features_din <= "0000100101111001";
        wait for Clk_period; 
        Features_din <= "1111101011010010";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "1111011001110000";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "1111110100110011";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000011101010";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000001001100000";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000001000111000";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000001001010101";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "1111011111011111";
        wait for Clk_period; 
        Features_din <= "0000000110010100";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111101111110111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000110011001001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000101011010110";
        wait for Clk_period; 
        Features_din <= "0000111011010010";
        wait for Clk_period; 
        Features_din <= "1111100000111100";
        wait for Clk_period; 
        Features_din <= "1111111000011110";
        wait for Clk_period; 
        Features_din <= "1111001100001100";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "1111100111110000";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000011110010";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000111010111";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000001011001";
        wait for Clk_period; 
        Features_din <= "1111100010100100";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101011011001";
        wait for Clk_period; 
        Features_din <= "0000001010000001";
        wait for Clk_period; 
        Features_din <= "0000001010000001";
        wait for Clk_period; 
        Features_din <= "0000001010000001";
        wait for Clk_period; 
        Features_din <= "0000001010000001";
        wait for Clk_period; 
        Features_din <= "0000001010000001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000100001011010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011010010001";
        wait for Clk_period; 
        Features_din <= "0000010100111011";
        wait for Clk_period; 
        Features_din <= "1111111000011111";
        wait for Clk_period; 
        Features_din <= "1111110001100011";
        wait for Clk_period; 
        Features_din <= "1111100011111010";
        wait for Clk_period; 
        Features_din <= "1111110100111100";
        wait for Clk_period; 
        Features_din <= "0000000100111001";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000010001011";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000001011010001";
        wait for Clk_period; 
        Features_din <= "0000000000101110";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000001011010100";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "1111100101101011";
        wait for Clk_period; 
        Features_din <= "0000001000111101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111100111110001";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001100110010100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111100001010";
        wait for Clk_period; 
        Features_din <= "0000001000001111";
        wait for Clk_period; 
        Features_din <= "1111001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "1111001000010111";
        wait for Clk_period; 
        Features_din <= "1111110101110111";
        wait for Clk_period; 
        Features_din <= "1111101000010000";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000101011101";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111011101011000";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110011101011";
        wait for Clk_period; 
        Features_din <= "0000001001011001";
        wait for Clk_period; 
        Features_din <= "0000001001011001";
        wait for Clk_period; 
        Features_din <= "0000001001011001";
        wait for Clk_period; 
        Features_din <= "0000001001011001";
        wait for Clk_period; 
        Features_din <= "0000001001011001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000101101001000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000111001100110";
        wait for Clk_period; 
        Features_din <= "0000011110011000";
        wait for Clk_period; 
        Features_din <= "1111011001101100";
        wait for Clk_period; 
        Features_din <= "0000000010101111";
        wait for Clk_period; 
        Features_din <= "1111100000010100";
        wait for Clk_period; 
        Features_din <= "1111111101110000";
        wait for Clk_period; 
        Features_din <= "1111111000000001";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000011100011";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "0000000010110011";
        wait for Clk_period; 
        Features_din <= "0000000101000001";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000110101011";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111011111010100";
        wait for Clk_period; 
        Features_din <= "0000000011111000";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111110000001001";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(3, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001000010010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001001000101";
        wait for Clk_period; 
        Features_din <= "0000111101001011";
        wait for Clk_period; 
        Features_din <= "1111110010111100";
        wait for Clk_period; 
        Features_din <= "0000001100000010";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "0000010010100100";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000010001110";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "0000001010001100";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "0000001100010101";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000010111000";
        wait for Clk_period; 
        Features_din <= "1111011111010100";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110000001001";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001100011111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000111101110011";
        wait for Clk_period; 
        Features_din <= "0000010010101011";
        wait for Clk_period; 
        Features_din <= "1111110101010110";
        wait for Clk_period; 
        Features_din <= "1111101011000001";
        wait for Clk_period; 
        Features_din <= "1111100011110111";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "1111101111001010";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000010101101";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000110101101";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "1111100000101100";
        wait for Clk_period; 
        Features_din <= "0000001001011000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101101111111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000100111100010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000111000111001";
        wait for Clk_period; 
        Features_din <= "0000101011110010";
        wait for Clk_period; 
        Features_din <= "1111011010111001";
        wait for Clk_period; 
        Features_din <= "1111111001010100";
        wait for Clk_period; 
        Features_din <= "1111001110011111";
        wait for Clk_period; 
        Features_din <= "1111111001110011";
        wait for Clk_period; 
        Features_din <= "0000000110101010";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000011011100";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000000011000000";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111011110101000";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110001010100";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000111001101111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000101010101100";
        wait for Clk_period; 
        Features_din <= "0000100110001000";
        wait for Clk_period; 
        Features_din <= "1111011001100111";
        wait for Clk_period; 
        Features_din <= "1111111101000111";
        wait for Clk_period; 
        Features_din <= "1111001001111101";
        wait for Clk_period; 
        Features_din <= "1111110000010001";
        wait for Clk_period; 
        Features_din <= "1111100010101100";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000011011011";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000001100000";
        wait for Clk_period; 
        Features_din <= "0000000010100000";
        wait for Clk_period; 
        Features_din <= "0000000011111010";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000100101010";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "1111011110000100";
        wait for Clk_period; 
        Features_din <= "0000000001111001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110010010100";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001000011000110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001000011100011";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "1110111111001001";
        wait for Clk_period; 
        Features_din <= "0000001100000011";
        wait for Clk_period; 
        Features_din <= "1111010010111110";
        wait for Clk_period; 
        Features_din <= "1111111110110011";
        wait for Clk_period; 
        Features_din <= "1111011010111000";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000011000001";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000000101011100";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000101111011";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "1111011101010010";
        wait for Clk_period; 
        Features_din <= "0000000010101100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110011110110";
        wait for Clk_period; 
        Features_din <= "0000001001011000";
        wait for Clk_period; 
        Features_din <= "0000001001011000";
        wait for Clk_period; 
        Features_din <= "0000001001011000";
        wait for Clk_period; 
        Features_din <= "0000001001011000";
        wait for Clk_period; 
        Features_din <= "0000001001011000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000110011110100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000000011001101";
        wait for Clk_period; 
        Features_din <= "0000100101110001";
        wait for Clk_period; 
        Features_din <= "1111110101001110";
        wait for Clk_period; 
        Features_din <= "1111110000100000";
        wait for Clk_period; 
        Features_din <= "1110110101001110";
        wait for Clk_period; 
        Features_din <= "1111101000011010";
        wait for Clk_period; 
        Features_din <= "1111111110000011";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000011100010";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000101101101";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "1111100000100100";
        wait for Clk_period; 
        Features_din <= "0000000101000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101110001010";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000101010000101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000100001000100";
        wait for Clk_period; 
        Features_din <= "0000011001101110";
        wait for Clk_period; 
        Features_din <= "1111011000010011";
        wait for Clk_period; 
        Features_din <= "1111110000011000";
        wait for Clk_period; 
        Features_din <= "1111010011010000";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000011011100";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000010000111";
        wait for Clk_period; 
        Features_din <= "0000000011010010";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000101001000";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000001000010101";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001100001100";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "1111100111110010";
        wait for Clk_period; 
        Features_din <= "0000001001000001";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111100101101010";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000110100101110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001001100000110";
        wait for Clk_period; 
        Features_din <= "0000000101010100";
        wait for Clk_period; 
        Features_din <= "1111010010101001";
        wait for Clk_period; 
        Features_din <= "0000010101000010";
        wait for Clk_period; 
        Features_din <= "1110111100100111";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "1111100001100001";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000011101011";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000010101001";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111011100110101";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110100110100";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001000001010010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111110010110110";
        wait for Clk_period; 
        Features_din <= "0000111101011011";
        wait for Clk_period; 
        Features_din <= "1111011001101111";
        wait for Clk_period; 
        Features_din <= "0000110000010001";
        wait for Clk_period; 
        Features_din <= "1111101101001000";
        wait for Clk_period; 
        Features_din <= "1111111001101111";
        wait for Clk_period; 
        Features_din <= "1111101100101101";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "0000000011001110";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "0000000000011010";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000110000010";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "1111011100110001";
        wait for Clk_period; 
        Features_din <= "0000000100000011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110100111100";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000001001010001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011110010011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010011011110";
        wait for Clk_period; 
        Features_din <= "0000100111000001";
        wait for Clk_period; 
        Features_din <= "1111011001101100";
        wait for Clk_period; 
        Features_din <= "1111111110111100";
        wait for Clk_period; 
        Features_din <= "1111011101010000";
        wait for Clk_period; 
        Features_din <= "0000000101011111";
        wait for Clk_period; 
        Features_din <= "0000001010101000";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000011011100";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000011000101";
        wait for Clk_period; 
        Features_din <= "0000000100001001";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000100000100";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "1111011111000011";
        wait for Clk_period; 
        Features_din <= "0000000010000100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110000100101";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000110011011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111011100010001";
        wait for Clk_period; 
        Features_din <= "0001001010010111";
        wait for Clk_period; 
        Features_din <= "1111001111100001";
        wait for Clk_period; 
        Features_din <= "0000100001001100";
        wait for Clk_period; 
        Features_din <= "0000011001101001";
        wait for Clk_period; 
        Features_din <= "0000001011111110";
        wait for Clk_period; 
        Features_din <= "1111101001100011";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000011000011";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "1111011100100101";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110101010111";
        wait for Clk_period; 
        Features_din <= "0000001001001110";
        wait for Clk_period; 
        Features_din <= "0000001001001110";
        wait for Clk_period; 
        Features_din <= "0000001001001110";
        wait for Clk_period; 
        Features_din <= "0000001001001110";
        wait for Clk_period; 
        Features_din <= "0000001001001110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001011111011110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000101010000110";
        wait for Clk_period; 
        Features_din <= "0000011101011110";
        wait for Clk_period; 
        Features_din <= "1110111110110101";
        wait for Clk_period; 
        Features_din <= "0000001010101101";
        wait for Clk_period; 
        Features_din <= "1111000001110011";
        wait for Clk_period; 
        Features_din <= "1111111010011110";
        wait for Clk_period; 
        Features_din <= "1111110011000011";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000011100001";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000101110100";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "1111100011010010";
        wait for Clk_period; 
        Features_din <= "0000000101000101";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111101010100000";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000010000101111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000110011101001";
        wait for Clk_period; 
        Features_din <= "0000010100001010";
        wait for Clk_period; 
        Features_din <= "1111100111000010";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "1111011111000111";
        wait for Clk_period; 
        Features_din <= "0000001000110110";
        wait for Clk_period; 
        Features_din <= "1111100010011100";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000011101111";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "1111011101100110";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110011001111";
        wait for Clk_period; 
        Features_din <= "0000001001011100";
        wait for Clk_period; 
        Features_din <= "0000001001011100";
        wait for Clk_period; 
        Features_din <= "0000001001011100";
        wait for Clk_period; 
        Features_din <= "0000001001011100";
        wait for Clk_period; 
        Features_din <= "0000001001011100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001100001000011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111110001111011";
        wait for Clk_period; 
        Features_din <= "0000100110010100";
        wait for Clk_period; 
        Features_din <= "1111010111010100";
        wait for Clk_period; 
        Features_din <= "0000000100100010";
        wait for Clk_period; 
        Features_din <= "1111110111000110";
        wait for Clk_period; 
        Features_din <= "1111011100100000";
        wait for Clk_period; 
        Features_din <= "1111100011101010";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000011100111";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "0000000000100101";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "1111011100010111";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111110101110111";
        wait for Clk_period; 
        Features_din <= "0000001001001010";
        wait for Clk_period; 
        Features_din <= "0000001001001010";
        wait for Clk_period; 
        Features_din <= "0000001001001010";
        wait for Clk_period; 
        Features_din <= "0000001001001010";
        wait for Clk_period; 
        Features_din <= "0000001001001010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001001000100000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001000110100100";
        wait for Clk_period; 
        Features_din <= "0000001001000101";
        wait for Clk_period; 
        Features_din <= "1111000001100101";
        wait for Clk_period; 
        Features_din <= "0000011111010111";
        wait for Clk_period; 
        Features_din <= "1111000010010001";
        wait for Clk_period; 
        Features_din <= "1111111100101111";
        wait for Clk_period; 
        Features_din <= "1111000101000100";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000011011110";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000000011000010";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "1111011011111010";
        wait for Clk_period; 
        Features_din <= "0000000000010010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110110111101";
        wait for Clk_period; 
        Features_din <= "0000001001000010";
        wait for Clk_period; 
        Features_din <= "0000001001000010";
        wait for Clk_period; 
        Features_din <= "0000001001000010";
        wait for Clk_period; 
        Features_din <= "0000001001000010";
        wait for Clk_period; 
        Features_din <= "0000001001000010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011100010010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001001011010011";
        wait for Clk_period; 
        Features_din <= "0000100010110001";
        wait for Clk_period; 
        Features_din <= "1111011110010100";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111010111011111";
        wait for Clk_period; 
        Features_din <= "0000001100010010";
        wait for Clk_period; 
        Features_din <= "1111011011011001";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000011100100";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000010100100";
        wait for Clk_period; 
        Features_din <= "0000000100010000";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000001011011";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000001001001111";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000001100010111";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111100001011000";
        wait for Clk_period; 
        Features_din <= "0000000100100110";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111101101000000";
        wait for Clk_period; 
        Features_din <= "0000001001111011";
        wait for Clk_period; 
        Features_din <= "0000001001111011";
        wait for Clk_period; 
        Features_din <= "0000001001111011";
        wait for Clk_period; 
        Features_din <= "0000001001111011";
        wait for Clk_period; 
        Features_din <= "0000001001111011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111110011011011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000110111001010";
        wait for Clk_period; 
        Features_din <= "1111111111100101";
        wait for Clk_period; 
        Features_din <= "1111111100101110";
        wait for Clk_period; 
        Features_din <= "1111011110000011";
        wait for Clk_period; 
        Features_din <= "1111010100111111";
        wait for Clk_period; 
        Features_din <= "1111011101100101";
        wait for Clk_period; 
        Features_din <= "0000100001101011";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000001011101";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000110111100";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "1111101000110011";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "1111100100101110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001000110001";
        wait for Clk_period; 
        Features_din <= "0000000101000111";
        wait for Clk_period; 
        Features_din <= "0000001100010111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001010011000111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111110111001011";
        wait for Clk_period; 
        Features_din <= "0000010010101100";
        wait for Clk_period; 
        Features_din <= "1111000101001010";
        wait for Clk_period; 
        Features_din <= "0000110010001001";
        wait for Clk_period; 
        Features_din <= "1111100010101100";
        wait for Clk_period; 
        Features_din <= "1111101100101110";
        wait for Clk_period; 
        Features_din <= "1111110011100100";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000000010001100";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000010111111";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "1111011101100100";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110011010011";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000001001011011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011100111000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000011010111101";
        wait for Clk_period; 
        Features_din <= "1111011111100101";
        wait for Clk_period; 
        Features_din <= "0000000100100011";
        wait for Clk_period; 
        Features_din <= "1111010011101000";
        wait for Clk_period; 
        Features_din <= "0000010111100101";
        wait for Clk_period; 
        Features_din <= "1111100101101100";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "1111011110000011";
        wait for Clk_period; 
        Features_din <= "0000000000010100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110010011000";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000001001100001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011100111111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000101001001000";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "1111110010011100";
        wait for Clk_period; 
        Features_din <= "1111110111100100";
        wait for Clk_period; 
        Features_din <= "1111100101011101";
        wait for Clk_period; 
        Features_din <= "1111110110010011";
        wait for Clk_period; 
        Features_din <= "0000000011010011";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000010111110";
        wait for Clk_period; 
        Features_din <= "0000000110000101";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000110111000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "1111100101100001";
        wait for Clk_period; 
        Features_din <= "0000000110000100";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111100111111011";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(3, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000100011001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111111111101000";
        wait for Clk_period; 
        Features_din <= "0000110001101000";
        wait for Clk_period; 
        Features_din <= "0001100010011111";
        wait for Clk_period; 
        Features_din <= "1111100001100011";
        wait for Clk_period; 
        Features_din <= "1111110001000101";
        wait for Clk_period; 
        Features_din <= "1111100010111100";
        wait for Clk_period; 
        Features_din <= "0000000011000111";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000000010001001";
        wait for Clk_period; 
        Features_din <= "0000000010110001";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000001010001";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "1111100001001101";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101101001111";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000001001111010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001010100000111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111110110011100";
        wait for Clk_period; 
        Features_din <= "0001000101001111";
        wait for Clk_period; 
        Features_din <= "1111011101100001";
        wait for Clk_period; 
        Features_din <= "0000100111100000";
        wait for Clk_period; 
        Features_din <= "1110110100111101";
        wait for Clk_period; 
        Features_din <= "0000010100010001";
        wait for Clk_period; 
        Features_din <= "1111010100000111";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000011100111";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000010100010";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000100010001";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "1111011111110011";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101111010101";
        wait for Clk_period; 
        Features_din <= "0000001001110001";
        wait for Clk_period; 
        Features_din <= "0000001001110001";
        wait for Clk_period; 
        Features_din <= "0000001001110001";
        wait for Clk_period; 
        Features_din <= "0000001001110001";
        wait for Clk_period; 
        Features_din <= "0000001001110001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000100100100111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0001000000100000";
        wait for Clk_period; 
        Features_din <= "1111110101111011";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "1111110001100110";
        wait for Clk_period; 
        Features_din <= "0000000110001011";
        wait for Clk_period; 
        Features_din <= "1111110111101010";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000011011100";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "0000000010110110";
        wait for Clk_period; 
        Features_din <= "0000000011111000";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000001011111110";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000001001111001";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000000000110001";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111100111111010";
        wait for Clk_period; 
        Features_din <= "0000000110000110";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "1111100101100010";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001101101110001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111010011110000";
        wait for Clk_period; 
        Features_din <= "0000010101000001";
        wait for Clk_period; 
        Features_din <= "1111011001101010";
        wait for Clk_period; 
        Features_din <= "1111111110101001";
        wait for Clk_period; 
        Features_din <= "1111011001110110";
        wait for Clk_period; 
        Features_din <= "0000000011011001";
        wait for Clk_period; 
        Features_din <= "0000001100010010";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000001100011";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000000011001100";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000110000001";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "1111100011101010";
        wait for Clk_period; 
        Features_din <= "0000000011100000";
        wait for Clk_period; 
        Features_din <= "0000000000011100";
        wait for Clk_period; 
        Features_din <= "1111101010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001101000111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000111010100111";
        wait for Clk_period; 
        Features_din <= "0000011001001010";
        wait for Clk_period; 
        Features_din <= "1111011101000101";
        wait for Clk_period; 
        Features_din <= "1111101110010111";
        wait for Clk_period; 
        Features_din <= "1111100000010001";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "0000010001111100";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000011100010";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001100111";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000001000101011";
        wait for Clk_period; 
        Features_din <= "0000000000110101";
        wait for Clk_period; 
        Features_din <= "0000000000010000";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000111110111";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000001010111010";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111100000011100";
        wait for Clk_period; 
        Features_din <= "0000000101001010";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111101110010111";
        wait for Clk_period; 
        Features_din <= "0000001001110110";
        wait for Clk_period; 
        Features_din <= "0000001001110110";
        wait for Clk_period; 
        Features_din <= "0000001001110110";
        wait for Clk_period; 
        Features_din <= "0000001001110110";
        wait for Clk_period; 
        Features_din <= "0000001001110110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000110010111110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000100110001101";
        wait for Clk_period; 
        Features_din <= "1111011111010000";
        wait for Clk_period; 
        Features_din <= "0000000010010011";
        wait for Clk_period; 
        Features_din <= "1111100011011001";
        wait for Clk_period; 
        Features_din <= "1111111100101011";
        wait for Clk_period; 
        Features_din <= "1111100101111111";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000000001111";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000010000110";
        wait for Clk_period; 
        Features_din <= "0000000010111100";
        wait for Clk_period; 
        Features_din <= "0000001000111100";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "1111011110001100";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110010000111";
        wait for Clk_period; 
        Features_din <= "0000001001100011";
        wait for Clk_period; 
        Features_din <= "0000001001100011";
        wait for Clk_period; 
        Features_din <= "0000001001100011";
        wait for Clk_period; 
        Features_din <= "0000001001100011";
        wait for Clk_period; 
        Features_din <= "0000001001100011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000000010101101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000100101010110";
        wait for Clk_period; 
        Features_din <= "0000001010100011";
        wait for Clk_period; 
        Features_din <= "1111100011111110";
        wait for Clk_period; 
        Features_din <= "1111101101001110";
        wait for Clk_period; 
        Features_din <= "1111100001110101";
        wait for Clk_period; 
        Features_din <= "1111101011101000";
        wait for Clk_period; 
        Features_din <= "0000001011011001";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000010111110";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "1111011110000110";
        wait for Clk_period; 
        Features_din <= "0000000000011001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110010010001";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000001001100010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000100100000101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000111010100100";
        wait for Clk_period; 
        Features_din <= "0000011110101100";
        wait for Clk_period; 
        Features_din <= "1111010101011010";
        wait for Clk_period; 
        Features_din <= "1111110101001111";
        wait for Clk_period; 
        Features_din <= "1111010100110100";
        wait for Clk_period; 
        Features_din <= "0000000101101110";
        wait for Clk_period; 
        Features_din <= "1111010011100111";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000011100011";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "0000000010101101";
        wait for Clk_period; 
        Features_din <= "0000000110000101";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000001001111101";
        wait for Clk_period; 
        Features_din <= "0000000001110111";
        wait for Clk_period; 
        Features_din <= "0000001010111101";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111100010011000";
        wait for Clk_period; 
        Features_din <= "0000001000100000";
        wait for Clk_period; 
        Features_din <= "0000000000001110";
        wait for Clk_period; 
        Features_din <= "1111101011101000";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000110011000001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000101000111011";
        wait for Clk_period; 
        Features_din <= "0000000100111110";
        wait for Clk_period; 
        Features_din <= "1111010000010001";
        wait for Clk_period; 
        Features_din <= "0000011110100000";
        wait for Clk_period; 
        Features_din <= "1111001100100011";
        wait for Clk_period; 
        Features_din <= "0000001100010110";
        wait for Clk_period; 
        Features_din <= "1111111011100000";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000010110100";
        wait for Clk_period; 
        Features_din <= "0000001011010111";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000001010111010";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000000010110101";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "1111100011011101";
        wait for Clk_period; 
        Features_din <= "0000000111110001";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "1111101010010010";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011000100011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011010011101";
        wait for Clk_period; 
        Features_din <= "0000011111010011";
        wait for Clk_period; 
        Features_din <= "1111101000101111";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "1111011010001011";
        wait for Clk_period; 
        Features_din <= "0000011100010101";
        wait for Clk_period; 
        Features_din <= "1111100111100001";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000011101010";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000000000100";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "1111011101110101";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110010110001";
        wait for Clk_period; 
        Features_din <= "0000001001011111";
        wait for Clk_period; 
        Features_din <= "0000001001011111";
        wait for Clk_period; 
        Features_din <= "0000001001011111";
        wait for Clk_period; 
        Features_din <= "0000001001011111";
        wait for Clk_period; 
        Features_din <= "0000001001011111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011011010001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000110011111011";
        wait for Clk_period; 
        Features_din <= "0000100000000010";
        wait for Clk_period; 
        Features_din <= "1111100100111000";
        wait for Clk_period; 
        Features_din <= "1111111011101100";
        wait for Clk_period; 
        Features_din <= "1111011110111101";
        wait for Clk_period; 
        Features_din <= "0000000101001111";
        wait for Clk_period; 
        Features_din <= "1111110110110111";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000011101011";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000010010010";
        wait for Clk_period; 
        Features_din <= "0000001010011100";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000111001011";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000001001110010";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001111000";
        wait for Clk_period; 
        Features_din <= "1111011110100011";
        wait for Clk_period; 
        Features_din <= "0000000110011010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110001011100";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011110011100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000111111001100";
        wait for Clk_period; 
        Features_din <= "0000011010100011";
        wait for Clk_period; 
        Features_din <= "1111100001000000";
        wait for Clk_period; 
        Features_din <= "1111101111100011";
        wait for Clk_period; 
        Features_din <= "1111100000010111";
        wait for Clk_period; 
        Features_din <= "1111110011111000";
        wait for Clk_period; 
        Features_din <= "1111101110001001";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000011110001";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000001101100";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000000110000110";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "1111100010010110";
        wait for Clk_period; 
        Features_din <= "0000001000111101";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101011101011";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001001110011110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011111000100";
        wait for Clk_period; 
        Features_din <= "0000100011010111";
        wait for Clk_period; 
        Features_din <= "1111001011110010";
        wait for Clk_period; 
        Features_din <= "0000100010111001";
        wait for Clk_period; 
        Features_din <= "1111001000010101";
        wait for Clk_period; 
        Features_din <= "0000010101001011";
        wait for Clk_period; 
        Features_din <= "1110111111100100";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000011100001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000011000010";
        wait for Clk_period; 
        Features_din <= "0000000011000000";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000000011101";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000111100011";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "1111011111010100";
        wait for Clk_period; 
        Features_din <= "0000000010100111";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111110000001001";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000100111101001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000110010001001";
        wait for Clk_period; 
        Features_din <= "0000011110000010";
        wait for Clk_period; 
        Features_din <= "1111101011100111";
        wait for Clk_period; 
        Features_din <= "1111111011110000";
        wait for Clk_period; 
        Features_din <= "1111000011100000";
        wait for Clk_period; 
        Features_din <= "0000000011110001";
        wait for Clk_period; 
        Features_din <= "1111101110001110";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000011110001";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001011010";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000000111111100";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000000111011010";
        wait for Clk_period; 
        Features_din <= "0000000001011111";
        wait for Clk_period; 
        Features_din <= "0000001011110000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "1111100000000000";
        wait for Clk_period; 
        Features_din <= "0000000100010100";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111101111000010";
        wait for Clk_period; 
        Features_din <= "0000001001110011";
        wait for Clk_period; 
        Features_din <= "0000001001110011";
        wait for Clk_period; 
        Features_din <= "0000001001110011";
        wait for Clk_period; 
        Features_din <= "0000001001110011";
        wait for Clk_period; 
        Features_din <= "0000001001110011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000100101000110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000101001010001";
        wait for Clk_period; 
        Features_din <= "0000010100101110";
        wait for Clk_period; 
        Features_din <= "1111011001001110";
        wait for Clk_period; 
        Features_din <= "0000100000001101";
        wait for Clk_period; 
        Features_din <= "1111011101101110";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "1111110001100110";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "0000000010100110";
        wait for Clk_period; 
        Features_din <= "0000000001001000";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "0000000001010011";
        wait for Clk_period; 
        Features_din <= "0000001100001101";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000001010000001";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "1111100011101000";
        wait for Clk_period; 
        Features_din <= "0000000100010100";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111101010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000101001110010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000110000111011";
        wait for Clk_period; 
        Features_din <= "0000001011101011";
        wait for Clk_period; 
        Features_din <= "1111101000100010";
        wait for Clk_period; 
        Features_din <= "1111110011000000";
        wait for Clk_period; 
        Features_din <= "1110111101000111";
        wait for Clk_period; 
        Features_din <= "1111111010110111";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000010001010";
        wait for Clk_period; 
        Features_din <= "0000000011000101";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000000100100";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000001100101";
        wait for Clk_period; 
        Features_din <= "1111011101110010";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110010111000";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000001001011110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000100000010011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000110110001000";
        wait for Clk_period; 
        Features_din <= "1111010101001111";
        wait for Clk_period; 
        Features_din <= "0000001100111000";
        wait for Clk_period; 
        Features_din <= "1111001101111011";
        wait for Clk_period; 
        Features_din <= "0000100101000101";
        wait for Clk_period; 
        Features_din <= "1111110001000100";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000011100001";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000010011100";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000010111111";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111100001100001";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000000010110";
        wait for Clk_period; 
        Features_din <= "1111101100110011";
        wait for Clk_period; 
        Features_din <= "0000001001111100";
        wait for Clk_period; 
        Features_din <= "0000001001111100";
        wait for Clk_period; 
        Features_din <= "0000001001111100";
        wait for Clk_period; 
        Features_din <= "0000001001111100";
        wait for Clk_period; 
        Features_din <= "0000001001111100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000010100010110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010111010100";
        wait for Clk_period; 
        Features_din <= "0000010010110100";
        wait for Clk_period; 
        Features_din <= "1111101101010100";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "1111100001001110";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "1111101010110111";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000010010101";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000001111101";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000000001101";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000001000000001";
        wait for Clk_period; 
        Features_din <= "0000000010000000";
        wait for Clk_period; 
        Features_din <= "0000000011011010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001111100";
        wait for Clk_period; 
        Features_din <= "1111011110011010";
        wait for Clk_period; 
        Features_din <= "0000000110101000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110001101100";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000001001100101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000111001001010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001000101010001";
        wait for Clk_period; 
        Features_din <= "0000000101111100";
        wait for Clk_period; 
        Features_din <= "1111010011000110";
        wait for Clk_period; 
        Features_din <= "1111011101100000";
        wait for Clk_period; 
        Features_din <= "1111011001011010";
        wait for Clk_period; 
        Features_din <= "0000000000101011";
        wait for Clk_period; 
        Features_din <= "1111100100101111";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000010111001";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000111100100";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000000001010";
        wait for Clk_period; 
        Features_din <= "0000000001001110";
        wait for Clk_period; 
        Features_din <= "0000001001001111";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000001010101010";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "1111011111010111";
        wait for Clk_period; 
        Features_din <= "0000000011010001";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111110000000011";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000001001101110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0001000100010010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001000010000111";
        wait for Clk_period; 
        Features_din <= "0000011111010110";
        wait for Clk_period; 
        Features_din <= "1111100100111101";
        wait for Clk_period; 
        Features_din <= "0000010001100001";
        wait for Clk_period; 
        Features_din <= "1111011011100011";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "1111011100111000";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "0000000111100000";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000110011110";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000000101010011";
        wait for Clk_period; 
        Features_din <= "0000001011100111";
        wait for Clk_period; 
        Features_din <= "0000000001001011";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "1111101010001101";
        wait for Clk_period; 
        Features_din <= "0000001000111010";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "1111100011100001";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000001010000100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(6, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "1111101110101100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "1111100010100100";
        wait for Clk_period; 
        Features_din <= "0000011001110100";
        wait for Clk_period; 
        Features_din <= "1111100001011011";
        wait for Clk_period; 
        Features_din <= "1111111001000001";
        wait for Clk_period; 
        Features_din <= "0001011000011011";
        wait for Clk_period; 
        Features_din <= "1111110100000011";
        wait for Clk_period; 
        Features_din <= "1111111101110010";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000010110111";
        wait for Clk_period; 
        Features_din <= "0000000011110000";
        wait for Clk_period; 
        Features_din <= "0000001100110010";
        wait for Clk_period; 
        Features_din <= "0000000000100001";
        wait for Clk_period; 
        Features_din <= "0000000000010101";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000100111011";
        wait for Clk_period; 
        Features_din <= "0000000010100001";
        wait for Clk_period; 
        Features_din <= "0000001000010010";
        wait for Clk_period; 
        Features_din <= "0000001011111101";
        wait for Clk_period; 
        Features_din <= "0000000000110100";
        wait for Clk_period; 
        Features_din <= "0000000001010100";
        wait for Clk_period; 
        Features_din <= "1111100011001010";
        wait for Clk_period; 
        Features_din <= "0000001010101000";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "1111101010101001";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000001010000011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000101001101100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010010000000";
        wait for Clk_period; 
        Features_din <= "0000101101100100";
        wait for Clk_period; 
        Features_din <= "1111001001000100";
        wait for Clk_period; 
        Features_din <= "0000001011111100";
        wait for Clk_period; 
        Features_din <= "1111010111111101";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "1111100011000110";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000011101001";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000010110010";
        wait for Clk_period; 
        Features_din <= "0000000000010011";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "0000000001100001";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000110111";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "1111011110100110";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110001010111";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000001001100111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011011110000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001000110101100";
        wait for Clk_period; 
        Features_din <= "0000010110001010";
        wait for Clk_period; 
        Features_din <= "1111011001011100";
        wait for Clk_period; 
        Features_din <= "1111110110001001";
        wait for Clk_period; 
        Features_din <= "1111010110011111";
        wait for Clk_period; 
        Features_din <= "1111111001001001";
        wait for Clk_period; 
        Features_din <= "0000001100110001";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000010101101";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000010001000";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000001001100";
        wait for Clk_period; 
        Features_din <= "0000000001101101";
        wait for Clk_period; 
        Features_din <= "0000000010000001";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111100001111001";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "1111101100010010";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000001001111110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000100000110111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011010001110";
        wait for Clk_period; 
        Features_din <= "0000101000111000";
        wait for Clk_period; 
        Features_din <= "1111011100110010";
        wait for Clk_period; 
        Features_din <= "1111111001001000";
        wait for Clk_period; 
        Features_din <= "1111011000000101";
        wait for Clk_period; 
        Features_din <= "0000000011100110";
        wait for Clk_period; 
        Features_din <= "1111110000111011";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000011011001";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000001110100";
        wait for Clk_period; 
        Features_din <= "0000000010110010";
        wait for Clk_period; 
        Features_din <= "0000000111111101";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000011111000";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000001001010101";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000001010010010";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "1111100100001010";
        wait for Clk_period; 
        Features_din <= "0000001000001100";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "1111101001011101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000101010001101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000110011101000";
        wait for Clk_period; 
        Features_din <= "0000010011110111";
        wait for Clk_period; 
        Features_din <= "1111100000101001";
        wait for Clk_period; 
        Features_din <= "0000000011011010";
        wait for Clk_period; 
        Features_din <= "1111001011001111";
        wait for Clk_period; 
        Features_din <= "1111110111110000";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "0000000001010111";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000000010010100";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "0000000001110101";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000010011000";
        wait for Clk_period; 
        Features_din <= "1111011111011111";
        wait for Clk_period; 
        Features_din <= "0000000000000011";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101111110101";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000110000110010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011010111000";
        wait for Clk_period; 
        Features_din <= "0000010100110100";
        wait for Clk_period; 
        Features_din <= "1111010011101011";
        wait for Clk_period; 
        Features_din <= "1111111001000011";
        wait for Clk_period; 
        Features_din <= "1111101011011110";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000111110111";
        wait for Clk_period; 
        Features_din <= "0000000000101100";
        wait for Clk_period; 
        Features_din <= "0000000011101111";
        wait for Clk_period; 
        Features_din <= "0000000000110110";
        wait for Clk_period; 
        Features_din <= "0000000010000011";
        wait for Clk_period; 
        Features_din <= "0000000100001101";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000000010010000";
        wait for Clk_period; 
        Features_din <= "0000000000101101";
        wait for Clk_period; 
        Features_din <= "0000000110110000";
        wait for Clk_period; 
        Features_din <= "0000000001110000";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000000000100111";
        wait for Clk_period; 
        Features_din <= "0000000001000000";
        wait for Clk_period; 
        Features_din <= "1111101001010110";
        wait for Clk_period; 
        Features_din <= "0000000100011100";
        wait for Clk_period; 
        Features_din <= "0000000010010110";
        wait for Clk_period; 
        Features_din <= "1111100100010000";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011010110011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001100010011100";
        wait for Clk_period; 
        Features_din <= "0000011101010100";
        wait for Clk_period; 
        Features_din <= "1111001101100000";
        wait for Clk_period; 
        Features_din <= "1111101111110101";
        wait for Clk_period; 
        Features_din <= "1111011001101100";
        wait for Clk_period; 
        Features_din <= "1111101101110011";
        wait for Clk_period; 
        Features_din <= "1111110010010100";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "0000001100011010";
        wait for Clk_period; 
        Features_din <= "0000000001001010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000001000101111";
        wait for Clk_period; 
        Features_din <= "0000000001101111";
        wait for Clk_period; 
        Features_din <= "0000000101000110";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "0000000010011010";
        wait for Clk_period; 
        Features_din <= "1111100001000001";
        wait for Clk_period; 
        Features_din <= "0000000101111010";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101101011111";
        wait for Clk_period; 
        Features_din <= "0000001001111001";
        wait for Clk_period; 
        Features_din <= "0000001001111001";
        wait for Clk_period; 
        Features_din <= "0000001001111001";
        wait for Clk_period; 
        Features_din <= "0000001001111001";
        wait for Clk_period; 
        Features_din <= "0000001001111001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000110011100011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000101000001111";
        wait for Clk_period; 
        Features_din <= "0000001011100001";
        wait for Clk_period; 
        Features_din <= "1111100111010100";
        wait for Clk_period; 
        Features_din <= "0000001001010111";
        wait for Clk_period; 
        Features_din <= "1111010101100110";
        wait for Clk_period; 
        Features_din <= "1111111100110001";
        wait for Clk_period; 
        Features_din <= "1111101001110101";
        wait for Clk_period; 
        Features_din <= "0000000000110011";
        wait for Clk_period; 
        Features_din <= "0000000011100000";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000010000101";
        wait for Clk_period; 
        Features_din <= "0000000011000111";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000000100000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111011";
        wait for Clk_period; 
        Features_din <= "0000000010100101";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000001010101";
        wait for Clk_period; 
        Features_din <= "1111011101000100";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110100010101";
        wait for Clk_period; 
        Features_din <= "0000001001010101";
        wait for Clk_period; 
        Features_din <= "0000001001010101";
        wait for Clk_period; 
        Features_din <= "0000001001010101";
        wait for Clk_period; 
        Features_din <= "0000001001010101";
        wait for Clk_period; 
        Features_din <= "0000001001010101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000110001111111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011110111101";
        wait for Clk_period; 
        Features_din <= "0000100010000100";
        wait for Clk_period; 
        Features_din <= "1111101011101110";
        wait for Clk_period; 
        Features_din <= "0000100100111000";
        wait for Clk_period; 
        Features_din <= "1111101000110011";
        wait for Clk_period; 
        Features_din <= "0000000111000111";
        wait for Clk_period; 
        Features_din <= "1111100001110001";
        wait for Clk_period; 
        Features_din <= "0000000001001001";
        wait for Clk_period; 
        Features_din <= "0000000001111010";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000001101011";
        wait for Clk_period; 
        Features_din <= "0000000010011001";
        wait for Clk_period; 
        Features_din <= "0000000101111001";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001011000";
        wait for Clk_period; 
        Features_din <= "0000001100010101";
        wait for Clk_period; 
        Features_din <= "0000000001110110";
        wait for Clk_period; 
        Features_din <= "0000001000010101";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000000001001101";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "1111100011111111";
        wait for Clk_period; 
        Features_din <= "0000000100100110";
        wait for Clk_period; 
        Features_din <= "0000000000000110";
        wait for Clk_period; 
        Features_din <= "1111101001101010";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000111100111100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000111011101010";
        wait for Clk_period; 
        Features_din <= "0000010111101111";
        wait for Clk_period; 
        Features_din <= "1111101001101000";
        wait for Clk_period; 
        Features_din <= "0000001011000001";
        wait for Clk_period; 
        Features_din <= "1111000110000100";
        wait for Clk_period; 
        Features_din <= "0000000000100011";
        wait for Clk_period; 
        Features_din <= "1111010000000101";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000011100000";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "0000000010101000";
        wait for Clk_period; 
        Features_din <= "0000000010011110";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000011011000";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000001010001010";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000001100000111";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000001101000";
        wait for Clk_period; 
        Features_din <= "1111100001101001";
        wait for Clk_period; 
        Features_din <= "0000000100010100";
        wait for Clk_period; 
        Features_din <= "0000000000001000";
        wait for Clk_period; 
        Features_din <= "1111101100101000";
        wait for Clk_period; 
        Features_din <= "0000001001111101";
        wait for Clk_period; 
        Features_din <= "0000001001111101";
        wait for Clk_period; 
        Features_din <= "0000001001111101";
        wait for Clk_period; 
        Features_din <= "0000001001111101";
        wait for Clk_period; 
        Features_din <= "0000001001111101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(6, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110000101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001000100110";
        wait for Clk_period; 
        Features_din <= "1111111110010100";
        wait for Clk_period; 
        Features_din <= "1111000111001011";
        wait for Clk_period; 
        Features_din <= "1111000011001100";
        wait for Clk_period; 
        Features_din <= "0000111011101100";
        wait for Clk_period; 
        Features_din <= "0000011110011110";
        wait for Clk_period; 
        Features_din <= "1111101100101110";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000010011011";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000010001101";
        wait for Clk_period; 
        Features_din <= "0000000100010110";
        wait for Clk_period; 
        Features_din <= "0000001100001010";
        wait for Clk_period; 
        Features_din <= "0000000000011011";
        wait for Clk_period; 
        Features_din <= "0000000001010010";
        wait for Clk_period; 
        Features_din <= "0000000000101010";
        wait for Clk_period; 
        Features_din <= "0000000101000000";
        wait for Clk_period; 
        Features_din <= "0000000010101010";
        wait for Clk_period; 
        Features_din <= "0000001001001000";
        wait for Clk_period; 
        Features_din <= "0000001011101100";
        wait for Clk_period; 
        Features_din <= "0000000000100010";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "1111100000101100";
        wait for Clk_period; 
        Features_din <= "0000001010110110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111101101111111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000111010001110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0001001101001111";
        wait for Clk_period; 
        Features_din <= "0000100111010010";
        wait for Clk_period; 
        Features_din <= "1111010110101101";
        wait for Clk_period; 
        Features_din <= "0000010011011111";
        wait for Clk_period; 
        Features_din <= "1111000011010000";
        wait for Clk_period; 
        Features_din <= "0000000110001110";
        wait for Clk_period; 
        Features_din <= "1110111111011101";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000011110100";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001011110";
        wait for Clk_period; 
        Features_din <= "0000000010011101";
        wait for Clk_period; 
        Features_din <= "0000000101101000";
        wait for Clk_period; 
        Features_din <= "0000000000111000";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "0000000001000100";
        wait for Clk_period; 
        Features_din <= "0000001000111001";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000001100000011";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "1111011111000011";
        wait for Clk_period; 
        Features_din <= "0000000011011000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110000100101";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "0000001001101011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000111000111110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000100011100111";
        wait for Clk_period; 
        Features_din <= "0000011001011110";
        wait for Clk_period; 
        Features_din <= "1111010100010001";
        wait for Clk_period; 
        Features_din <= "1111111001011110";
        wait for Clk_period; 
        Features_din <= "1111010011010100";
        wait for Clk_period; 
        Features_din <= "1111110110110100";
        wait for Clk_period; 
        Features_din <= "1111101010001100";
        wait for Clk_period; 
        Features_din <= "0000000000111101";
        wait for Clk_period; 
        Features_din <= "0000000011101001";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001101010";
        wait for Clk_period; 
        Features_din <= "0000000010100011";
        wait for Clk_period; 
        Features_din <= "0000000000101001";
        wait for Clk_period; 
        Features_din <= "0000000000101111";
        wait for Clk_period; 
        Features_din <= "0000000000000010";
        wait for Clk_period; 
        Features_din <= "0000000001000101";
        wait for Clk_period; 
        Features_din <= "0000000011001000";
        wait for Clk_period; 
        Features_din <= "0000000001110010";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000111100";
        wait for Clk_period; 
        Features_din <= "0000000001101001";
        wait for Clk_period; 
        Features_din <= "1111011011111001";
        wait for Clk_period; 
        Features_din <= "0000000000011110";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "1111110111000000";
        wait for Clk_period; 
        Features_din <= "0000001001000001";
        wait for Clk_period; 
        Features_din <= "0000001001000001";
        wait for Clk_period; 
        Features_din <= "0000001001000001";
        wait for Clk_period; 
        Features_din <= "0000001001000001";
        wait for Clk_period; 
        Features_din <= "0000001001000001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000011110111101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000011101101011";
        wait for Clk_period; 
        Features_din <= "0000011010110010";
        wait for Clk_period; 
        Features_din <= "1111101000000100";
        wait for Clk_period; 
        Features_din <= "1111110110101000";
        wait for Clk_period; 
        Features_din <= "1111100000011111";
        wait for Clk_period; 
        Features_din <= "0000000011110101";
        wait for Clk_period; 
        Features_din <= "1111110101001000";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000011101101";
        wait for Clk_period; 
        Features_din <= "0000000000111111";
        wait for Clk_period; 
        Features_din <= "0000000001100100";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000000000001011";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000100011010";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000110111100";
        wait for Clk_period; 
        Features_din <= "0000000001110001";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000000000111110";
        wait for Clk_period; 
        Features_din <= "0000000001101110";
        wait for Clk_period; 
        Features_din <= "1111100101100010";
        wait for Clk_period; 
        Features_din <= "0000000110101101";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111100111111010";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000111011011001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        Features_din <= "0000101100111110";
        wait for Clk_period; 
        Features_din <= "1111100001000101";
        wait for Clk_period; 
        Features_din <= "0000011100110101";
        wait for Clk_period; 
        Features_din <= "1111011010111100";
        wait for Clk_period; 
        Features_din <= "0000001000010101";
        wait for Clk_period; 
        Features_din <= "1111100011011011";
        wait for Clk_period; 
        Features_din <= "0000000001000010";
        wait for Clk_period; 
        Features_din <= "0000000011011011";
        wait for Clk_period; 
        Features_din <= "0000000001000110";
        wait for Clk_period; 
        Features_din <= "0000000001111011";
        wait for Clk_period; 
        Features_din <= "0000000010111011";
        wait for Clk_period; 
        Features_din <= "0000000000000111";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "0000000011010101";
        wait for Clk_period; 
        Features_din <= "0000000000111001";
        wait for Clk_period; 
        Features_din <= "0000000110101011";
        wait for Clk_period; 
        Features_din <= "0000000001111111";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000000000110010";
        wait for Clk_period; 
        Features_din <= "0000000001010110";
        wait for Clk_period; 
        Features_din <= "1111100101111100";
        wait for Clk_period; 
        Features_din <= "0000000011010110";
        wait for Clk_period; 
        Features_din <= "0000000000100110";
        wait for Clk_period; 
        Features_din <= "1111100111011111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(7, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000101011110101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000110111000100";
        wait for Clk_period; 
        Features_din <= "0000011100000010";
        wait for Clk_period; 
        Features_din <= "1111100010111000";
        wait for Clk_period; 
        Features_din <= "0000000010010111";
        wait for Clk_period; 
        Features_din <= "1111010100011111";
        wait for Clk_period; 
        Features_din <= "1111110101111100";
        wait for Clk_period; 
        Features_din <= "1111110011000000";
        wait for Clk_period; 
        Features_din <= "0000000001000111";
        wait for Clk_period; 
        Features_din <= "0000000010110000";
        wait for Clk_period; 
        Features_din <= "0000000001000001";
        wait for Clk_period; 
        Features_din <= "0000000001110011";
        wait for Clk_period; 
        Features_din <= "0000000010111111";
        wait for Clk_period; 
        Features_din <= "0000000011010100";
        wait for Clk_period; 
        Features_din <= "0000000000110000";
        wait for Clk_period; 
        Features_din <= "0000000000001001";
        wait for Clk_period; 
        Features_din <= "0000000001000011";
        wait for Clk_period; 
        Features_din <= "0000000100001101";
        wait for Clk_period; 
        Features_din <= "0000000010000010";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000000000111010";
        wait for Clk_period; 
        Features_din <= "0000000001100110";
        wait for Clk_period; 
        Features_din <= "1111100000101011";
        wait for Clk_period; 
        Features_din <= "0000000001100010";
        wait for Clk_period; 
        Features_din <= "0000000000000001";
        wait for Clk_period; 
        Features_din <= "1111101110000000";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000001001110111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000000000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
            wait;
    end process;
end;
