

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.types.all;

entity image_test is
    generic(TREE_RAM_BITS: positive := 13;
            NUM_CLASSES:   positive := 7;
            NUM_FEATURES:  positive := 255);
end image_test;

architecture behavior of image_test is
    
    component image
        generic(TREE_RAM_BITS: positive;
                NUM_CLASSES:   positive;
                NUM_FEATURES:  positive);
        port(-- Control signals
             Clk:   in std_logic;
             Reset: in std_logic;
             
             -- Inputs for the nodes reception (trees)
             Load_trees: in std_logic;
             Valid_node: in std_logic;
             Addr:       in std_logic_vector(TREE_RAM_BITS - 1  downto 0);
             Trees_din:  in std_logic_vector(31 downto 0);
             
             -- Inputs for the features reception (pixels)
             Load_features: in std_logic;
             Valid_feature: in std_logic;
             Features_din:  in std_logic_vector(15 downto 0);
             Last_feature:  in std_logic;
             
             -- Output signals
             --     Finish:     finish (also 'ready') signal
             --     Dout:       the selected class
             --     Greater:    the value of the selected class prediction
             --     Curr_state: the current state
             Finish:     out std_logic;
             Dout:       out std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);
             greater:    out std_logic_vector(31 downto 0);
             curr_state: out std_logic_vector(2 downto 0));
    end component;
    
    component counter is
        generic(BITS: natural);
        port(Clk:   in  std_logic;
             Reset: in  std_logic;
             Count: in  std_logic;
             Dout:  out std_logic_vector (BITS - 1 downto 0));
    end component;
    
    -- Inputs
    signal Clk:           std_logic := '0';
    signal Reset:         std_logic := '0';
    signal Load_trees:    std_logic := '0';
    signal Valid_node:    std_logic := '0';
    signal Addr:          std_logic_vector(TREE_RAM_BITS - 1 downto
                                           0) := (others => '0');
    signal Trees_din:     std_logic_vector(31 downto 0) := (others => '0');
    signal Load_features: std_logic := '0';
    signal Valid_feature: std_logic := '0';
    signal Features_din:  std_logic_vector(15 downto 0) := (others => '0');
    signal last_feature:  std_logic := '0';
    
    -- Outputs
    signal Finish:     std_logic;
    signal Dout:       std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);
    signal greater:    std_logic_vector(31 downto 0);
    signal curr_state: std_logic_vector(2 downto 0);
    
    -- Clock period definition
    constant Clk_period : time := 10 ns;
    
    -- Counter signals
    signal pc_count, hc_count: std_logic := '0';
    signal pixels, hits: std_logic_vector(15 downto 0) := (others => '0');
    
    -- Label signal
    signal class_label: std_logic_vector(log_2(NUM_CLASSES) - 1 downto 0);

begin
    
    -- Instantiate the Unit Under Test (UUT)
    uut: image
        generic map(TREE_RAM_BITS => TREE_RAM_BITS,
                    NUM_CLASSES   => NUM_CLASSES,
                    NUM_FEATURES  => NUM_FEATURES)
        port map(Clk           => Clk,
                 Reset         => Reset,
                 Load_trees    => Load_trees,
                 Valid_node    => Valid_node,
                 Addr          => Addr,
                 Trees_din     => Trees_din,
                 Load_features => Load_features,
                 Valid_feature => Valid_feature,
                 Features_din  => Features_din,
                 Last_feature  => Last_feature,
                 Finish        => Finish,
                 Dout          => Dout,
                 greater       => greater,
                 curr_state    => curr_state);
    
    -- To count the pixels
    pixel_counter: counter
        generic map(BITS => 16)
        port map(Clk   => Clk, 
                 Reset => Reset,
                 Count => pc_count,
                 Dout  => pixels);
    
    -- To count the hits
    hit_counter: counter
        generic map(BITS => 16)
        port map(Clk   => Clk, 
                 Reset => Reset,
                 Count => hc_count,
                 Dout  => hits);
    
    -- Clock process definition
    Clk_process: process
    begin
        Clk <= '0';
        wait for Clk_period/2;
        Clk <= '1';
        wait for Clk_period/2;
    end process;
    
    -- Stimulus process
    stim_proc: process
    begin
        
        Reset <= '1';
        
        -- hold reset state for 100 ns.
        wait for 100 ns;
        
        Reset <= '0';
        
        wait for Clk_period*10;
        


        
        -- LOAD TREES
        -----------------------------------------------------------------------
        
        -- Load and valid trees flags
        Load_trees <= '1';
        Valid_node <= '1';

        -- Class  0
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"0a0a3664";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"1e079e38";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"9e06511c";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"5f0c6f10";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"150abb08";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"63000204";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"ffc2011d";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"ff51011d";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"0701ae04";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"01c6011d";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"ff8f011d";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"d9095c08";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"0a097204";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"ff71011d";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"0027011d";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"0280011d";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"15059110";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"0a070208";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"0b00dc04";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"01a3011d";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"ff62011d";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"d9047704";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"ff89011d";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"02fb011d";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"d6052508";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"49015604";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"ff95011d";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"0391011d";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"ff71011d";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"2a050518";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"5f08bf10";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"28074708";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"55001504";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"0027011d";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"ff52011d";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"03010904";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"01c6011d";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"ff81011d";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"16046f04";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"0332011d";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"ff78011d";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"5100f108";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"0c015c04";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"013c011d";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"ff61011d";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"16087c08";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"4e045a04";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"0059011d";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"03e2011d";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"ff8f011d";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"52022f24";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"69005d08";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"0b012104";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"ff7a011d";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"0027011d";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"7202350c";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"980a9808";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"25006a04";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"0154011d";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"0421011d";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"0071011d";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"0604d508";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"0300cd04";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"0027011d";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"ff7d011d";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"1f00d604";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"00b2011d";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"036c011d";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"23072504";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"ff54011d";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"0154011d";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"95060f48";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"0a08ea2c";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"0609eb20";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"5f0b0010";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"9e086e08";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"5f054b04";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"ff560249";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"ff850249";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"0b013904";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"01400249";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"ff7e0249";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"1d070908";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"50005004";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"00340249";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"ff770249";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"3b017304";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"019e0249";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"00190249";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"68020308";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"a5049704";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"008b0249";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"01d60249";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"ff6f0249";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"0e03ff0c";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"e7027d04";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"ff580249";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"48012004";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"017b0249";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"ff9f0249";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"a706c00c";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"3b022608";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"6803ee04";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"01bf0249";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"00150249";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"fffa0249";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"ff870249";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"b405c530";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"4e07ca1c";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"28070b10";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"d109eb08";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"1d07d504";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"ff590249";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"00370249";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"0a097204";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"ffa90249";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"00fc0249";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"37026508";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"1c02e304";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"01af0249";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"002e0249";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"ff8c0249";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"0a043008";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"1e0b1304";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"ff670249";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"00ca0249";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"51010004";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"ff800249";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"f9005104";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"ff940249";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"019e0249";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"4901770c";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"c100f408";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"06070a04";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"000f0249";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"00ff0249";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"ff620249";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"52030e10";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"25008b08";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"2807c404";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"ff790249";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"01170249";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"09007504";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"ff8c0249";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"01b00249";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"ff7b0249";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"9505ac54";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"3b00fc2c";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"49031d14";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"0608c90c";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"5f088a04";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"ff59038d";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"2900df04";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"00b2038d";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"0005038d";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"31028c04";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"ffa5038d";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"010e038d";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"6d034908";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"db0b5504";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"ff69038d";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"002d038d";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"5a054f08";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"7202b904";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"0143038d";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"ffb7038d";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"02005504";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"00a0038d";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"ff73038d";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"6300000c";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"96012f08";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"2201b004";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"0202038d";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"001c038d";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"ff6f038d";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"3700430c";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"2e008a08";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"5701a204";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"014f038d";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"ff97038d";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"ff5f038d";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"2807eb08";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"6d0d1f04";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"ff5a038d";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"0006038d";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"5a012004";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"00c3038d";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"ff5e038d";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"4e053a24";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"1d06d014";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"2807930c";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"9e083f04";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"ff59038d";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"0a028904";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"ff85038d";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"00cb038d";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"91054b04";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"0007038d";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"012e038d";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"6802c00c";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"0b06e608";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"c8005f04";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"004e038d";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"015d038d";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"ff9e038d";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"ff86038d";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"0900c20c";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"24101304";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"ff5e038d";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"0b06e604";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"00cb038d";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"fffd038d";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"ac035a10";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"77015708";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"9d004804";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"012d038d";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"ff97038d";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"37004a04";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"00c6038d";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"ff6e038d";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"4900ea08";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"d3000004";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"0029038d";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"ff8a038d";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"26040804";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"0135038d";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"ff97038d";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"6d060e48";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"9e07a12c";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"1508d41c";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"66005410";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"37014908";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"d1069704";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"fff204a9";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"01a304a9";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"d601a404";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"003204a9";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"ff6204a9";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"1d0ed808";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"63000904";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"ffba04a9";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"ff5e04a9";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"006204a9";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"0e03b804";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"ff6b04a9";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"a0005208";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"f1003904";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"007104a9";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"ff8e04a9";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"013304a9";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"ee082714";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"06034208";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"fb038004";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"ff7f04a9";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"002d04a9";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"5e031608";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"73012604";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"005a04a9";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"011704a9";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"fff504a9";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"1e089804";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"ff6104a9";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"002f04a9";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"15023720";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"950a4f10";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"5f091308";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"46002604";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"fffc04a9";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"ff5c04a9";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"83000004";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"00d304a9";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"ff6e04a9";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"5a097c0c";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"9e036a04";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"ffdc04a9";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"79044404";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"004904a9";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"00f504a9";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"ff7e04a9";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"0e033710";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"3b009408";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"0d020504";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"00c804a9";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"001604a9";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"db0a8f04";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"ff6304a9";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"007604a9";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"c107d810";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"fe033408";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"49016f04";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"fffa04a9";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"00fe04a9";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"62005004";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"006c04a9";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"ff7504a9";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"dc00c104";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"002204a9";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"ff6e04a9";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"7604903c";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"0e04b320";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"6600480c";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"37015d08";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"7d020704";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"ffaa05bd";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"012105bd";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"ff6c05bd";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"1e08c30c";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"3c0c8c08";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"5d10a304";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"ff5f05bd";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"001705bd";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"000805bd";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"52003804";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"009305bd";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"ff9305bd";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"ea03bc14";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"59021910";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"ac01bc08";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"0a063804";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"ff8b05bd";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"005205bd";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"cd018404";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"002205bd";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"00fe05bd";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"ff7005bd";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"67000504";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"006005bd";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"ff5f05bd";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"0a044624";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"0b01ff14";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"5200e10c";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"7a02c308";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"0301ed04";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"011b05bd";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"fff505bd";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"ff9c05bd";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"00014f04";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"003405bd";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"ff6f05bd";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"0609eb08";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"9008eb04";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"ff5f05bd";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"003e05bd";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"840e2904";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"ff9c05bd";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"00be05bd";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"0e034f10";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"cc00f808";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"d107b704";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"ffa305bd";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"00d405bd";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"71009504";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"001505bd";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"ff6905bd";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"1605dc10";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"c8002a08";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"b302c304";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"009505bd";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"ff7105bd";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"09005c04";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"ffa105bd";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"00dd05bd";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"c7014a08";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"24032c04";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"ffa005bd";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"00c005bd";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"ff6d05bd";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"76049058";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"9e03e528";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"3b00ab10";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"0a04b304";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"ff7206f1";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"c9039804";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"ff9106f1";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"b2035304";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"003406f1";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"010006f1";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"6600480c";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"8b010908";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"43009404";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"00c606f1";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"ffeb06f1";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"ff7406f1";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"5f0d0508";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"8b0bf104";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"ff6006f1";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"ffb806f1";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"001606f1";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"0a07201c";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"1505a50c";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"17000a08";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"09028204";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"ff9806f1";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"009d06f1";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"ff6106f1";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"cb02e608";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"5a02c104";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"00c606f1";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"ffa606f1";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"b5005a04";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"fff306f1";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"ff7a06f1";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"25009c08";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"54004e04";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"ffff06f1";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"ff8606f1";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"0c030e08";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"2e030f04";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"00df06f1";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"ffe106f1";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"ffcb06f1";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"0a02df14";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"0b01600c";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"00012608";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"ee07e504";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"00ea06f1";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"001e06f1";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"ff8006f1";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"490ac604";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"ff6206f1";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"005506f1";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"59020918";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"4900ea08";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"86000004";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"000d06f1";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"ff7506f1";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"0e034f08";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"cc00f804";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"009906f1";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"ff9606f1";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"2d0a2604";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"00c706f1";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"ff9206f1";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"1d05ce08";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"890c3b04";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"ff6806f1";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"ffee06f1";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"c502c808";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"db035604";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"ffa106f1";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"00b006f1";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"1b017604";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"ff7806f1";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"fffb06f1";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"76049040";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"0e04b324";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"66008b14";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"cc01f410";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"c5016b08";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"f000b904";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"015307fd";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"005707fd";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"9e05e004";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"ff8707fd";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"003707fd";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"ff6f07fd";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"a4003a04";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"001607fd";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"2a0c9508";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"5d10a304";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"ff6207fd";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"000807fd";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"000d07fd";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"ea03bc14";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"59021910";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"6d037308";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"0b03ab04";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"ffa007fd";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"001907fd";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"7301ef04";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"ffeb07fd";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"00c907fd";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"ff7e07fd";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"06081104";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"ff6507fd";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"002c07fd";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"15023724";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"2a06a814";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"0a076608";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"06089504";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"ff6507fd";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"000907fd";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"ac084508";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"b6019d04";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"ff8a07fd";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"ffe107fd";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"008d07fd";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"3b016908";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"9d07f704";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"00be07fd";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"ffa907fd";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"3b042504";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"ff7b07fd";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"ffee07fd";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"0c031d14";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"2d093110";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"0e033708";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"ce016c04";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"006a07fd";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"ff8007fd";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"09007504";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"ff9b07fd";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"00b707fd";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"ff8407fd";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"23074e08";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"68004404";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"002507fd";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"ff6e07fd";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"5a01ce04";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"009e07fd";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"ffc707fd";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"6d053840";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"3b011d1c";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"2a036008";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"760b7904";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"ff6c091d";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"fff3091d";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"00010e0c";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"0901fc04";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"ff9f091d";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"6b039d04";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"0026091d";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"00d8091d";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"1d07d504";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"ff80091d";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"005c091d";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"2806db14";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"9e097b0c";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"790b7e08";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"47001a04";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"ffe4091d";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"ff64091d";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"0002091d";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"ea060e04";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"0065091d";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"ffa1091d";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"76049008";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"ba000a04";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"003a091d";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"ff6e091d";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"55029204";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"00f9091d";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"ffb1091d";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"0a054524";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"0b029f18";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"cd027b08";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"cf00e104";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"0028091d";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"ff77091d";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"9d043208";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"9e036a04";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"ffeb091d";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"00b6091d";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"1f0da104";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"ff93091d";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"0047091d";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"06096108";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"90083604";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"ff66091d";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"0049091d";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"0065091d";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"2602d020";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"15020010";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"ad013b08";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"4e060904";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"ffc5091d";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"0093091d";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"e4062d04";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"ff75091d";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"0036091d";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"3d04d508";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"65001104";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"ffd4091d";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"00ae091d";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"fa00e704";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"fffe091d";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"ff9e091d";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"2309e808";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"fd022704";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"ff71091d";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"0033091d";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"0094091d";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"1e046040";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"5f06b324";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"0608c918";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"66008b0c";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"67008d04";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"00960a39";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"72001a04";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"001c0a39";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"ff760a39";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"6d0e2608";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"0a0b7704";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"ff650a39";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"ffd70a39";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"00050a39";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"3b007e04";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"00820a39";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"05029904";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"ff970a39";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"ffee0a39";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"24038a0c";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"3b00a304";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"002d0a39";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"2e000104";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"fff80a39";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"ff6b0a39";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"15022e04";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"ff890a39";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"2601d808";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"73037604";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"000c0a39";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"00bb0a39";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"ffad0a39";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"ac034828";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"4e07ca14";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"3b01600c";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"b3022f04";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"ff830a39";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"2f028404";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"00890a39";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"ffae0a39";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"4e070904";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"ff680a39";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"ffde0a39";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"eb039710";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"c904b908";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"b406c904";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"ff9e0a39";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"00630a39";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"5a023304";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"00d40a39";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"002a0a39";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"ff8a0a39";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"0901e614";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"7303ae0c";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"2d013504";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"00210a39";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"cc000004";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"ffdc0a39";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"ff740a39";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"06020f04";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"ffce0a39";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"007a0a39";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"65001d08";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"df001804";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"007e0a39";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"ff890a39";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"2d0a2608";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"69004804";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"fff30a39";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"00a80a39";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"ffb20a39";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"1e04493c";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"5f06b328";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"0608c91c";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"66008b10";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"2106b208";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"9107e804";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"ff7d0b45";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"ffe40b45";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"cc02ac04";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"00f50b45";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"ffb00b45";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"0a0b7708";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"74096704";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"ff660b45";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"ffc30b45";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"ffe00b45";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"ce009b04";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"006f0b45";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"ae023304";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"ffa30b45";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"ffea0b45";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"15022e04";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"ff7b0b45";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"26019b08";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"73030304";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"ffc90b45";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"00a50b45";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"2d00e104";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"ff840b45";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"00050b45";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"ac028620";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"1d07fb14";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"59009710";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"3806da08";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"5c026c04";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"ff850b45";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"ffed0b45";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"d3006b04";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"007a0b45";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"00000b45";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"ff6b0b45";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"0202d604";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"ffaf0b45";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"5a023f04";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"00990b45";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"00240b45";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"0a057c14";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"0b04c710";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"25027508";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"4c030604";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"ffec0b45";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"ff840b45";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"06029704";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"ffae0b45";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"008d0b45";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"ff7a0b45";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"ef023210";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"5b044f08";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"0901e604";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"001f0b45";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"00a40b45";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"1e077004";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"ff9d0b45";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"00500b45";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"7606e104";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"ff860b45";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"00540b45";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"0a070258";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"4e06ce24";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"63001c0c";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"e2030808";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"40007e04";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"000a0c51";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"ff7a0c51";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"00c70c51";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"1e079e0c";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"3a000404";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"ffe70c51";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"0609eb04";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"ff660c51";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"ffd50c51";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"0b016b08";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"c7022704";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"00630c51";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"ffcb0c51";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"ff8a0c51";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"0301ed18";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"c7019010";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"0e044a08";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"d8000c04";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"00530c51";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"ffa90c51";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"0b03ab04";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"00ad0c51";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"00120c51";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"3808e704";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"ff930c51";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"003c0c51";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"760a4310";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"15061a08";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"a3049104";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"ff6d0c51";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"ffdb0c51";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"49051704";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"ffeb0c51";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"001c0c51";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"2a025604";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"ffa70c51";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"e00a6704";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"007a0c51";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"00040c51";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"26023420";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"e5035410";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"3d03b80c";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"980a9808";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"65001304";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"ffe60c51";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"00a10c51";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"ffdc0c51";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"ffe90c51";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"23074e08";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"38076904";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"ff940c51";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"00170c51";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"82038704";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"ffee0c51";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"008b0c51";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"2306eb08";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"0e05a104";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"ff6f0c51";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"00240c51";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"a0001604";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"ffe00c51";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"007e0c51";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"1e044930";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"5f06b31c";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"0608c914";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"66008b08";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"2106b204";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"ff940d35";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"00750d35";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"5f065108";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"d10a8e04";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"ff680d35";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"ffd50d35";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"ffde0d35";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"07027a04";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"00510d35";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"ffb20d35";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"15022e04";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"ff880d35";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"b601c308";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"0d029404";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"00990d35";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"fff00d35";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"d500c904";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"ff900d35";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"001e0d35";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"4e04e614";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"2807c40c";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"1d074104";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"ff700d35";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"00005404";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"00670d35";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"ffdf0d35";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"62011f04";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"00800d35";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"00020d35";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"0a059518";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"b405c50c";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"ac052804";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"ff7f0d35";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"0b020904";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"00480d35";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"ffaa0d35";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"4900da04";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"ffa50d35";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"7002ae04";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"00810d35";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"ffd70d35";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"59028a0c";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"8803b808";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"0900f704";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"ffee0d35";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"009a0d35";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"ffc40d35";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"be007a04";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"ff8e0d35";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"71042d04";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"005e0d35";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"00140d35";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"1e04492c";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"5e018e1c";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"0b02f114";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"24036b08";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"a2035c04";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"ff970e11";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"000c0e11";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"1b01e308";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"02018904";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"00370e11";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"00d50e11";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"00260e11";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"2d00cd04";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"000a0e11";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"ff790e11";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"0a0b210c";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"8d001f04";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"ffda0e11";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"2d000004";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"ffd50e11";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"ff680e11";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"000a0e11";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"0e03a214";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"71024a0c";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"2304e304";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"ffa20e11";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"db07b604";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"00120e11";
		wait for Clk_period;
		Addr <=  "0001101101001";
		Trees_din <= x"00750e11";
		wait for Clk_period;
		Addr <=  "0001101101010";
		Trees_din <= x"d10a5904";
		wait for Clk_period;
		Addr <=  "0001101101011";
		Trees_din <= x"ff730e11";
		wait for Clk_period;
		Addr <=  "0001101101100";
		Trees_din <= x"fff10e11";
		wait for Clk_period;
		Addr <=  "0001101101101";
		Trees_din <= x"2a060318";
		wait for Clk_period;
		Addr <=  "0001101101110";
		Trees_din <= x"2d020e0c";
		wait for Clk_period;
		Addr <=  "0001101101111";
		Trees_din <= x"0e050004";
		wait for Clk_period;
		Addr <=  "0001101110000";
		Trees_din <= x"ffd30e11";
		wait for Clk_period;
		Addr <=  "0001101110001";
		Trees_din <= x"2e032504";
		wait for Clk_period;
		Addr <=  "0001101110010";
		Trees_din <= x"00820e11";
		wait for Clk_period;
		Addr <=  "0001101110011";
		Trees_din <= x"00110e11";
		wait for Clk_period;
		Addr <=  "0001101110100";
		Trees_din <= x"9e083f04";
		wait for Clk_period;
		Addr <=  "0001101110101";
		Trees_din <= x"ff820e11";
		wait for Clk_period;
		Addr <=  "0001101110110";
		Trees_din <= x"d40af904";
		wait for Clk_period;
		Addr <=  "0001101110111";
		Trees_din <= x"ffb40e11";
		wait for Clk_period;
		Addr <=  "0001101111000";
		Trees_din <= x"00480e11";
		wait for Clk_period;
		Addr <=  "0001101111001";
		Trees_din <= x"5902010c";
		wait for Clk_period;
		Addr <=  "0001101111010";
		Trees_din <= x"8803b808";
		wait for Clk_period;
		Addr <=  "0001101111011";
		Trees_din <= x"30050c04";
		wait for Clk_period;
		Addr <=  "0001101111100";
		Trees_din <= x"009f0e11";
		wait for Clk_period;
		Addr <=  "0001101111101";
		Trees_din <= x"00310e11";
		wait for Clk_period;
		Addr <=  "0001101111110";
		Trees_din <= x"ffdb0e11";
		wait for Clk_period;
		Addr <=  "0001101111111";
		Trees_din <= x"be005704";
		wait for Clk_period;
		Addr <=  "0001110000000";
		Trees_din <= x"ffac0e11";
		wait for Clk_period;
		Addr <=  "0001110000001";
		Trees_din <= x"1d086204";
		wait for Clk_period;
		Addr <=  "0001110000010";
		Trees_din <= x"001c0e11";
		wait for Clk_period;
		Addr <=  "0001110000011";
		Trees_din <= x"007b0e11";
		wait for Clk_period;
		Addr <=  "0001110000100";
		Trees_din <= x"0a068330";
		wait for Clk_period;
		Addr <=  "0001110000101";
		Trees_din <= x"0e05ec14";
		wait for Clk_period;
		Addr <=  "0001110000110";
		Trees_din <= x"0300430c";
		wait for Clk_period;
		Addr <=  "0001110000111";
		Trees_din <= x"67006d04";
		wait for Clk_period;
		Addr <=  "0001110001000";
		Trees_din <= x"00780ecd";
		wait for Clk_period;
		Addr <=  "0001110001001";
		Trees_din <= x"3e01ee04";
		wait for Clk_period;
		Addr <=  "0001110001010";
		Trees_din <= x"ffe10ecd";
		wait for Clk_period;
		Addr <=  "0001110001011";
		Trees_din <= x"ff840ecd";
		wait for Clk_period;
		Addr <=  "0001110001100";
		Trees_din <= x"8b000804";
		wait for Clk_period;
		Addr <=  "0001110001101";
		Trees_din <= x"fffb0ecd";
		wait for Clk_period;
		Addr <=  "0001110001110";
		Trees_din <= x"ff6a0ecd";
		wait for Clk_period;
		Addr <=  "0001110001111";
		Trees_din <= x"49025908";
		wait for Clk_period;
		Addr <=  "0001110010000";
		Trees_din <= x"0e131404";
		wait for Clk_period;
		Addr <=  "0001110010001";
		Trees_din <= x"ff790ecd";
		wait for Clk_period;
		Addr <=  "0001110010010";
		Trees_din <= x"00000ecd";
		wait for Clk_period;
		Addr <=  "0001110010011";
		Trees_din <= x"9d04d00c";
		wait for Clk_period;
		Addr <=  "0001110010100";
		Trees_din <= x"0601ae04";
		wait for Clk_period;
		Addr <=  "0001110010101";
		Trees_din <= x"fff60ecd";
		wait for Clk_period;
		Addr <=  "0001110010110";
		Trees_din <= x"9e036a04";
		wait for Clk_period;
		Addr <=  "0001110010111";
		Trees_din <= x"001f0ecd";
		wait for Clk_period;
		Addr <=  "0001110011000";
		Trees_din <= x"008d0ecd";
		wait for Clk_period;
		Addr <=  "0001110011001";
		Trees_din <= x"06063504";
		wait for Clk_period;
		Addr <=  "0001110011010";
		Trees_din <= x"ff9e0ecd";
		wait for Clk_period;
		Addr <=  "0001110011011";
		Trees_din <= x"00150ecd";
		wait for Clk_period;
		Addr <=  "0001110011100";
		Trees_din <= x"26024e20";
		wait for Clk_period;
		Addr <=  "0001110011101";
		Trees_din <= x"e5035414";
		wait for Clk_period;
		Addr <=  "0001110011110";
		Trees_din <= x"c8002608";
		wait for Clk_period;
		Addr <=  "0001110011111";
		Trees_din <= x"52004704";
		wait for Clk_period;
		Addr <=  "0001110100000";
		Trees_din <= x"00490ecd";
		wait for Clk_period;
		Addr <=  "0001110100001";
		Trees_din <= x"ffbb0ecd";
		wait for Clk_period;
		Addr <=  "0001110100010";
		Trees_din <= x"0900f704";
		wait for Clk_period;
		Addr <=  "0001110100011";
		Trees_din <= x"ffe70ecd";
		wait for Clk_period;
		Addr <=  "0001110100100";
		Trees_din <= x"a1084c04";
		wait for Clk_period;
		Addr <=  "0001110100101";
		Trees_din <= x"00970ecd";
		wait for Clk_period;
		Addr <=  "0001110100110";
		Trees_din <= x"fff40ecd";
		wait for Clk_period;
		Addr <=  "0001110100111";
		Trees_din <= x"0604b104";
		wait for Clk_period;
		Addr <=  "0001110101000";
		Trees_din <= x"ffa90ecd";
		wait for Clk_period;
		Addr <=  "0001110101001";
		Trees_din <= x"2f01fa04";
		wait for Clk_period;
		Addr <=  "0001110101010";
		Trees_din <= x"00690ecd";
		wait for Clk_period;
		Addr <=  "0001110101011";
		Trees_din <= x"ffda0ecd";
		wait for Clk_period;
		Addr <=  "0001110101100";
		Trees_din <= x"2306eb08";
		wait for Clk_period;
		Addr <=  "0001110101101";
		Trees_din <= x"0a0e2c04";
		wait for Clk_period;
		Addr <=  "0001110101110";
		Trees_din <= x"ff7a0ecd";
		wait for Clk_period;
		Addr <=  "0001110101111";
		Trees_din <= x"fffa0ecd";
		wait for Clk_period;
		Addr <=  "0001110110000";
		Trees_din <= x"bf00aa04";
		wait for Clk_period;
		Addr <=  "0001110110001";
		Trees_din <= x"fffc0ecd";
		wait for Clk_period;
		Addr <=  "0001110110010";
		Trees_din <= x"00660ecd";
		wait for Clk_period;
		Addr <=  "0001110110011";
		Trees_din <= x"1e044924";
		wait for Clk_period;
		Addr <=  "0001110110100";
		Trees_din <= x"63001c0c";
		wait for Clk_period;
		Addr <=  "0001110110101";
		Trees_din <= x"9a020b08";
		wait for Clk_period;
		Addr <=  "0001110110110";
		Trees_din <= x"fb03de04";
		wait for Clk_period;
		Addr <=  "0001110110111";
		Trees_din <= x"00120f81";
		wait for Clk_period;
		Addr <=  "0001110111000";
		Trees_din <= x"00aa0f81";
		wait for Clk_period;
		Addr <=  "0001110111001";
		Trees_din <= x"ffaf0f81";
		wait for Clk_period;
		Addr <=  "0001110111010";
		Trees_din <= x"0606d510";
		wait for Clk_period;
		Addr <=  "0001110111011";
		Trees_din <= x"380b0908";
		wait for Clk_period;
		Addr <=  "0001110111100";
		Trees_din <= x"3b004c04";
		wait for Clk_period;
		Addr <=  "0001110111101";
		Trees_din <= x"ffd70f81";
		wait for Clk_period;
		Addr <=  "0001110111110";
		Trees_din <= x"ff6d0f81";
		wait for Clk_period;
		Addr <=  "0001110111111";
		Trees_din <= x"6c023604";
		wait for Clk_period;
		Addr <=  "0001111000000";
		Trees_din <= x"002f0f81";
		wait for Clk_period;
		Addr <=  "0001111000001";
		Trees_din <= x"ffb50f81";
		wait for Clk_period;
		Addr <=  "0001111000010";
		Trees_din <= x"d905ce04";
		wait for Clk_period;
		Addr <=  "0001111000011";
		Trees_din <= x"ffa60f81";
		wait for Clk_period;
		Addr <=  "0001111000100";
		Trees_din <= x"00540f81";
		wait for Clk_period;
		Addr <=  "0001111000101";
		Trees_din <= x"4e04e60c";
		wait for Clk_period;
		Addr <=  "0001111000110";
		Trees_din <= x"2807c408";
		wait for Clk_period;
		Addr <=  "0001111000111";
		Trees_din <= x"1d074104";
		wait for Clk_period;
		Addr <=  "0001111001000";
		Trees_din <= x"ff7a0f81";
		wait for Clk_period;
		Addr <=  "0001111001001";
		Trees_din <= x"002a0f81";
		wait for Clk_period;
		Addr <=  "0001111001010";
		Trees_din <= x"004d0f81";
		wait for Clk_period;
		Addr <=  "0001111001011";
		Trees_din <= x"2a058118";
		wait for Clk_period;
		Addr <=  "0001111001100";
		Trees_din <= x"57026710";
		wait for Clk_period;
		Addr <=  "0001111001101";
		Trees_din <= x"27067108";
		wait for Clk_period;
		Addr <=  "0001111001110";
		Trees_din <= x"53044c04";
		wait for Clk_period;
		Addr <=  "0001111001111";
		Trees_din <= x"fffc0f81";
		wait for Clk_period;
		Addr <=  "0001111010000";
		Trees_din <= x"007a0f81";
		wait for Clk_period;
		Addr <=  "0001111010001";
		Trees_din <= x"0a078304";
		wait for Clk_period;
		Addr <=  "0001111010010";
		Trees_din <= x"ffae0f81";
		wait for Clk_period;
		Addr <=  "0001111010011";
		Trees_din <= x"00060f81";
		wait for Clk_period;
		Addr <=  "0001111010100";
		Trees_din <= x"6c016504";
		wait for Clk_period;
		Addr <=  "0001111010101";
		Trees_din <= x"fff90f81";
		wait for Clk_period;
		Addr <=  "0001111010110";
		Trees_din <= x"ff960f81";
		wait for Clk_period;
		Addr <=  "0001111010111";
		Trees_din <= x"8803180c";
		wait for Clk_period;
		Addr <=  "0001111011000";
		Trees_din <= x"c8002604";
		wait for Clk_period;
		Addr <=  "0001111011001";
		Trees_din <= x"fff80f81";
		wait for Clk_period;
		Addr <=  "0001111011010";
		Trees_din <= x"3d02e604";
		wait for Clk_period;
		Addr <=  "0001111011011";
		Trees_din <= x"00920f81";
		wait for Clk_period;
		Addr <=  "0001111011100";
		Trees_din <= x"000c0f81";
		wait for Clk_period;
		Addr <=  "0001111011101";
		Trees_din <= x"0e063504";
		wait for Clk_period;
		Addr <=  "0001111011110";
		Trees_din <= x"ffab0f81";
		wait for Clk_period;
		Addr <=  "0001111011111";
		Trees_din <= x"00540f81";
		wait for Clk_period;
		Addr <=  "0001111100000";
		Trees_din <= x"0a068330";
		wait for Clk_period;
		Addr <=  "0001111100001";
		Trees_din <= x"e5019e1c";
		wait for Clk_period;
		Addr <=  "0001111100010";
		Trees_din <= x"49021c08";
		wait for Clk_period;
		Addr <=  "0001111100011";
		Trees_din <= x"18002c04";
		wait for Clk_period;
		Addr <=  "0001111100100";
		Trees_din <= x"ffea103d";
		wait for Clk_period;
		Addr <=  "0001111100101";
		Trees_din <= x"ff87103d";
		wait for Clk_period;
		Addr <=  "0001111100110";
		Trees_din <= x"38052c08";
		wait for Clk_period;
		Addr <=  "0001111100111";
		Trees_din <= x"47008204";
		wait for Clk_period;
		Addr <=  "0001111101000";
		Trees_din <= x"0024103d";
		wait for Clk_period;
		Addr <=  "0001111101001";
		Trees_din <= x"ffa4103d";
		wait for Clk_period;
		Addr <=  "0001111101010";
		Trees_din <= x"57026708";
		wait for Clk_period;
		Addr <=  "0001111101011";
		Trees_din <= x"59018604";
		wait for Clk_period;
		Addr <=  "0001111101100";
		Trees_din <= x"0093103d";
		wait for Clk_period;
		Addr <=  "0001111101101";
		Trees_din <= x"0017103d";
		wait for Clk_period;
		Addr <=  "0001111101110";
		Trees_din <= x"fffc103d";
		wait for Clk_period;
		Addr <=  "0001111101111";
		Trees_din <= x"0e065f08";
		wait for Clk_period;
		Addr <=  "0001111110000";
		Trees_din <= x"df003104";
		wait for Clk_period;
		Addr <=  "0001111110001";
		Trees_din <= x"fff7103d";
		wait for Clk_period;
		Addr <=  "0001111110010";
		Trees_din <= x"ff6b103d";
		wait for Clk_period;
		Addr <=  "0001111110011";
		Trees_din <= x"49026404";
		wait for Clk_period;
		Addr <=  "0001111110100";
		Trees_din <= x"ff98103d";
		wait for Clk_period;
		Addr <=  "0001111110101";
		Trees_din <= x"2a06a804";
		wait for Clk_period;
		Addr <=  "0001111110110";
		Trees_din <= x"ffed103d";
		wait for Clk_period;
		Addr <=  "0001111110111";
		Trees_din <= x"0052103d";
		wait for Clk_period;
		Addr <=  "0001111111000";
		Trees_din <= x"3d01cc24";
		wait for Clk_period;
		Addr <=  "0001111111001";
		Trees_din <= x"cd011908";
		wait for Clk_period;
		Addr <=  "0001111111010";
		Trees_din <= x"47015a04";
		wait for Clk_period;
		Addr <=  "0001111111011";
		Trees_din <= x"003d103d";
		wait for Clk_period;
		Addr <=  "0001111111100";
		Trees_din <= x"ffaf103d";
		wait for Clk_period;
		Addr <=  "0001111111101";
		Trees_din <= x"5b029f0c";
		wait for Clk_period;
		Addr <=  "0001111111110";
		Trees_din <= x"aa010e04";
		wait for Clk_period;
		Addr <=  "0001111111111";
		Trees_din <= x"0015103d";
		wait for Clk_period;
		Addr <=  "0010000000000";
		Trees_din <= x"6803ee04";
		wait for Clk_period;
		Addr <=  "0010000000001";
		Trees_din <= x"0098103d";
		wait for Clk_period;
		Addr <=  "0010000000010";
		Trees_din <= x"002e103d";
		wait for Clk_period;
		Addr <=  "0010000000011";
		Trees_din <= x"23074e08";
		wait for Clk_period;
		Addr <=  "0010000000100";
		Trees_din <= x"eb00f604";
		wait for Clk_period;
		Addr <=  "0010000000101";
		Trees_din <= x"ffbd103d";
		wait for Clk_period;
		Addr <=  "0010000000110";
		Trees_din <= x"0013103d";
		wait for Clk_period;
		Addr <=  "0010000000111";
		Trees_din <= x"d107b704";
		wait for Clk_period;
		Addr <=  "0010000001000";
		Trees_din <= x"0018103d";
		wait for Clk_period;
		Addr <=  "0010000001001";
		Trees_din <= x"005b103d";
		wait for Clk_period;
		Addr <=  "0010000001010";
		Trees_din <= x"0e063504";
		wait for Clk_period;
		Addr <=  "0010000001011";
		Trees_din <= x"ff90103d";
		wait for Clk_period;
		Addr <=  "0010000001100";
		Trees_din <= x"9105a704";
		wait for Clk_period;
		Addr <=  "0010000001101";
		Trees_din <= x"ffed103d";
		wait for Clk_period;
		Addr <=  "0010000001110";
		Trees_din <= x"005b103d";
		wait for Clk_period;
		Addr <=  "0010000001111";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0010000010000";
		Trees_din <= x"0a06832c";
		wait for Clk_period;
		Addr <=  "0010000010001";
		Trees_din <= x"e5019e1c";
		wait for Clk_period;
		Addr <=  "0010000010010";
		Trees_din <= x"49021c08";
		wait for Clk_period;
		Addr <=  "0010000010011";
		Trees_din <= x"ec10a604";
		wait for Clk_period;
		Addr <=  "0010000010100";
		Trees_din <= x"ff8f10e5";
		wait for Clk_period;
		Addr <=  "0010000010101";
		Trees_din <= x"ffe510e5";
		wait for Clk_period;
		Addr <=  "0010000010110";
		Trees_din <= x"38052c08";
		wait for Clk_period;
		Addr <=  "0010000010111";
		Trees_din <= x"4700c204";
		wait for Clk_period;
		Addr <=  "0010000011000";
		Trees_din <= x"001a10e5";
		wait for Clk_period;
		Addr <=  "0010000011001";
		Trees_din <= x"ffab10e5";
		wait for Clk_period;
		Addr <=  "0010000011010";
		Trees_din <= x"0001fa08";
		wait for Clk_period;
		Addr <=  "0010000011011";
		Trees_din <= x"70027004";
		wait for Clk_period;
		Addr <=  "0010000011100";
		Trees_din <= x"008510e5";
		wait for Clk_period;
		Addr <=  "0010000011101";
		Trees_din <= x"000910e5";
		wait for Clk_period;
		Addr <=  "0010000011110";
		Trees_din <= x"ffe610e5";
		wait for Clk_period;
		Addr <=  "0010000011111";
		Trees_din <= x"28080f08";
		wait for Clk_period;
		Addr <=  "0010000100000";
		Trees_din <= x"240a7204";
		wait for Clk_period;
		Addr <=  "0010000100001";
		Trees_din <= x"ff7110e5";
		wait for Clk_period;
		Addr <=  "0010000100010";
		Trees_din <= x"fff910e5";
		wait for Clk_period;
		Addr <=  "0010000100011";
		Trees_din <= x"ad019204";
		wait for Clk_period;
		Addr <=  "0010000100100";
		Trees_din <= x"003d10e5";
		wait for Clk_period;
		Addr <=  "0010000100101";
		Trees_din <= x"ffb210e5";
		wait for Clk_period;
		Addr <=  "0010000100110";
		Trees_din <= x"c8002d08";
		wait for Clk_period;
		Addr <=  "0010000100111";
		Trees_din <= x"62011f04";
		wait for Clk_period;
		Addr <=  "0010000101000";
		Trees_din <= x"002f10e5";
		wait for Clk_period;
		Addr <=  "0010000101001";
		Trees_din <= x"ff9210e5";
		wait for Clk_period;
		Addr <=  "0010000101010";
		Trees_din <= x"37023e10";
		wait for Clk_period;
		Addr <=  "0010000101011";
		Trees_din <= x"d1021604";
		wait for Clk_period;
		Addr <=  "0010000101100";
		Trees_din <= x"ffe210e5";
		wait for Clk_period;
		Addr <=  "0010000101101";
		Trees_din <= x"62034708";
		wait for Clk_period;
		Addr <=  "0010000101110";
		Trees_din <= x"66041204";
		wait for Clk_period;
		Addr <=  "0010000101111";
		Trees_din <= x"009210e5";
		wait for Clk_period;
		Addr <=  "0010000110000";
		Trees_din <= x"002710e5";
		wait for Clk_period;
		Addr <=  "0010000110001";
		Trees_din <= x"000410e5";
		wait for Clk_period;
		Addr <=  "0010000110010";
		Trees_din <= x"23059408";
		wait for Clk_period;
		Addr <=  "0010000110011";
		Trees_din <= x"cb02a904";
		wait for Clk_period;
		Addr <=  "0010000110100";
		Trees_din <= x"000610e5";
		wait for Clk_period;
		Addr <=  "0010000110101";
		Trees_din <= x"ff9d10e5";
		wait for Clk_period;
		Addr <=  "0010000110110";
		Trees_din <= x"a2027404";
		wait for Clk_period;
		Addr <=  "0010000110111";
		Trees_din <= x"fff410e5";
		wait for Clk_period;
		Addr <=  "0010000111000";
		Trees_din <= x"006210e5";
		wait for Clk_period;
		Addr <=  "0010000111001";
		Trees_din <= x"2a067e2c";
		wait for Clk_period;
		Addr <=  "0010000111010";
		Trees_din <= x"e5019e18";
		wait for Clk_period;
		Addr <=  "0010000111011";
		Trees_din <= x"1504860c";
		wait for Clk_period;
		Addr <=  "0010000111100";
		Trees_din <= x"240b3208";
		wait for Clk_period;
		Addr <=  "0010000111101";
		Trees_din <= x"79047c04";
		wait for Clk_period;
		Addr <=  "0010000111110";
		Trees_din <= x"ff8f1189";
		wait for Clk_period;
		Addr <=  "0010000111111";
		Trees_din <= x"fff81189";
		wait for Clk_period;
		Addr <=  "0010001000000";
		Trees_din <= x"00241189";
		wait for Clk_period;
		Addr <=  "0010001000001";
		Trees_din <= x"38044f04";
		wait for Clk_period;
		Addr <=  "0010001000010";
		Trees_din <= x"ffec1189";
		wait for Clk_period;
		Addr <=  "0010001000011";
		Trees_din <= x"c4020904";
		wait for Clk_period;
		Addr <=  "0010001000100";
		Trees_din <= x"007b1189";
		wait for Clk_period;
		Addr <=  "0010001000101";
		Trees_din <= x"001e1189";
		wait for Clk_period;
		Addr <=  "0010001000110";
		Trees_din <= x"0606c10c";
		wait for Clk_period;
		Addr <=  "0010001000111";
		Trees_din <= x"d909c908";
		wait for Clk_period;
		Addr <=  "0010001001000";
		Trees_din <= x"0a089404";
		wait for Clk_period;
		Addr <=  "0010001001001";
		Trees_din <= x"ff6f1189";
		wait for Clk_period;
		Addr <=  "0010001001010";
		Trees_din <= x"ffcf1189";
		wait for Clk_period;
		Addr <=  "0010001001011";
		Trees_din <= x"fff61189";
		wait for Clk_period;
		Addr <=  "0010001001100";
		Trees_din <= x"6d054b04";
		wait for Clk_period;
		Addr <=  "0010001001101";
		Trees_din <= x"ffca1189";
		wait for Clk_period;
		Addr <=  "0010001001110";
		Trees_din <= x"00321189";
		wait for Clk_period;
		Addr <=  "0010001001111";
		Trees_din <= x"0e03a210";
		wait for Clk_period;
		Addr <=  "0010001010000";
		Trees_din <= x"71024a08";
		wait for Clk_period;
		Addr <=  "0010001010001";
		Trees_din <= x"8f01c104";
		wait for Clk_period;
		Addr <=  "0010001010010";
		Trees_din <= x"ffe91189";
		wait for Clk_period;
		Addr <=  "0010001010011";
		Trees_din <= x"00571189";
		wait for Clk_period;
		Addr <=  "0010001010100";
		Trees_din <= x"be008e04";
		wait for Clk_period;
		Addr <=  "0010001010101";
		Trees_din <= x"ff8f1189";
		wait for Clk_period;
		Addr <=  "0010001010110";
		Trees_din <= x"ffe01189";
		wait for Clk_period;
		Addr <=  "0010001010111";
		Trees_din <= x"59020110";
		wait for Clk_period;
		Addr <=  "0010001011000";
		Trees_din <= x"ee09f00c";
		wait for Clk_period;
		Addr <=  "0010001011001";
		Trees_din <= x"99000804";
		wait for Clk_period;
		Addr <=  "0010001011010";
		Trees_din <= x"00061189";
		wait for Clk_period;
		Addr <=  "0010001011011";
		Trees_din <= x"72027d04";
		wait for Clk_period;
		Addr <=  "0010001011100";
		Trees_din <= x"00921189";
		wait for Clk_period;
		Addr <=  "0010001011101";
		Trees_din <= x"00241189";
		wait for Clk_period;
		Addr <=  "0010001011110";
		Trees_din <= x"fff81189";
		wait for Clk_period;
		Addr <=  "0010001011111";
		Trees_din <= x"e0009f04";
		wait for Clk_period;
		Addr <=  "0010001100000";
		Trees_din <= x"ffb11189";
		wait for Clk_period;
		Addr <=  "0010001100001";
		Trees_din <= x"00351189";
		wait for Clk_period;
		Addr <=  "0010001100010";
		Trees_din <= x"0a05fe1c";
		wait for Clk_period;
		Addr <=  "0010001100011";
		Trees_din <= x"3805ab0c";
		wait for Clk_period;
		Addr <=  "0010001100100";
		Trees_din <= x"03001d04";
		wait for Clk_period;
		Addr <=  "0010001100101";
		Trees_din <= x"00031205";
		wait for Clk_period;
		Addr <=  "0010001100110";
		Trees_din <= x"d40af904";
		wait for Clk_period;
		Addr <=  "0010001100111";
		Trees_din <= x"ff751205";
		wait for Clk_period;
		Addr <=  "0010001101000";
		Trees_din <= x"ffd61205";
		wait for Clk_period;
		Addr <=  "0010001101001";
		Trees_din <= x"5a010c08";
		wait for Clk_period;
		Addr <=  "0010001101010";
		Trees_din <= x"00016804";
		wait for Clk_period;
		Addr <=  "0010001101011";
		Trees_din <= x"00721205";
		wait for Clk_period;
		Addr <=  "0010001101100";
		Trees_din <= x"ffea1205";
		wait for Clk_period;
		Addr <=  "0010001101101";
		Trees_din <= x"00003404";
		wait for Clk_period;
		Addr <=  "0010001101110";
		Trees_din <= x"001d1205";
		wait for Clk_period;
		Addr <=  "0010001101111";
		Trees_din <= x"ff981205";
		wait for Clk_period;
		Addr <=  "0010001110000";
		Trees_din <= x"2303ed08";
		wait for Clk_period;
		Addr <=  "0010001110001";
		Trees_din <= x"6e012004";
		wait for Clk_period;
		Addr <=  "0010001110010";
		Trees_din <= x"00271205";
		wait for Clk_period;
		Addr <=  "0010001110011";
		Trees_din <= x"ff9d1205";
		wait for Clk_period;
		Addr <=  "0010001110100";
		Trees_din <= x"5b026e10";
		wait for Clk_period;
		Addr <=  "0010001110101";
		Trees_din <= x"0901e604";
		wait for Clk_period;
		Addr <=  "0010001110110";
		Trees_din <= x"fff91205";
		wait for Clk_period;
		Addr <=  "0010001110111";
		Trees_din <= x"d3031908";
		wait for Clk_period;
		Addr <=  "0010001111000";
		Trees_din <= x"3d021f04";
		wait for Clk_period;
		Addr <=  "0010001111001";
		Trees_din <= x"008d1205";
		wait for Clk_period;
		Addr <=  "0010001111010";
		Trees_din <= x"001d1205";
		wait for Clk_period;
		Addr <=  "0010001111011";
		Trees_din <= x"000d1205";
		wait for Clk_period;
		Addr <=  "0010001111100";
		Trees_din <= x"59017b08";
		wait for Clk_period;
		Addr <=  "0010001111101";
		Trees_din <= x"0d01b404";
		wait for Clk_period;
		Addr <=  "0010001111110";
		Trees_din <= x"00571205";
		wait for Clk_period;
		Addr <=  "0010001111111";
		Trees_din <= x"fffb1205";
		wait for Clk_period;
		Addr <=  "0010010000000";
		Trees_din <= x"ffb81205";
		wait for Clk_period;
		Addr <=  "0010010000001";
		Trees_din <= x"1e044914";
		wait for Clk_period;
		Addr <=  "0010010000010";
		Trees_din <= x"63001c08";
		wait for Clk_period;
		Addr <=  "0010010000011";
		Trees_din <= x"80010d04";
		wait for Clk_period;
		Addr <=  "0010010000100";
		Trees_din <= x"00561279";
		wait for Clk_period;
		Addr <=  "0010010000101";
		Trees_din <= x"fff21279";
		wait for Clk_period;
		Addr <=  "0010010000110";
		Trees_din <= x"0606d508";
		wait for Clk_period;
		Addr <=  "0010010000111";
		Trees_din <= x"380b0904";
		wait for Clk_period;
		Addr <=  "0010010001000";
		Trees_din <= x"ff7c1279";
		wait for Clk_period;
		Addr <=  "0010010001001";
		Trees_din <= x"fff41279";
		wait for Clk_period;
		Addr <=  "0010010001010";
		Trees_din <= x"00001279";
		wait for Clk_period;
		Addr <=  "0010010001011";
		Trees_din <= x"ac02860c";
		wait for Clk_period;
		Addr <=  "0010010001100";
		Trees_din <= x"1d07fb08";
		wait for Clk_period;
		Addr <=  "0010010001101";
		Trees_din <= x"0e04d404";
		wait for Clk_period;
		Addr <=  "0010010001110";
		Trees_din <= x"ff931279";
		wait for Clk_period;
		Addr <=  "0010010001111";
		Trees_din <= x"ffef1279";
		wait for Clk_period;
		Addr <=  "0010010010000";
		Trees_din <= x"002f1279";
		wait for Clk_period;
		Addr <=  "0010010010001";
		Trees_din <= x"73019e08";
		wait for Clk_period;
		Addr <=  "0010010010010";
		Trees_din <= x"0604d504";
		wait for Clk_period;
		Addr <=  "0010010010011";
		Trees_din <= x"ffb31279";
		wait for Clk_period;
		Addr <=  "0010010010100";
		Trees_din <= x"000d1279";
		wait for Clk_period;
		Addr <=  "0010010010101";
		Trees_din <= x"72028410";
		wait for Clk_period;
		Addr <=  "0010010010110";
		Trees_din <= x"8802da08";
		wait for Clk_period;
		Addr <=  "0010010010111";
		Trees_din <= x"2802d604";
		wait for Clk_period;
		Addr <=  "0010010011000";
		Trees_din <= x"00171279";
		wait for Clk_period;
		Addr <=  "0010010011001";
		Trees_din <= x"00831279";
		wait for Clk_period;
		Addr <=  "0010010011010";
		Trees_din <= x"ca006804";
		wait for Clk_period;
		Addr <=  "0010010011011";
		Trees_din <= x"ffdd1279";
		wait for Clk_period;
		Addr <=  "0010010011100";
		Trees_din <= x"00391279";
		wait for Clk_period;
		Addr <=  "0010010011101";
		Trees_din <= x"ffda1279";
		wait for Clk_period;
		Addr <=  "0010010011110";
		Trees_din <= x"15042318";
		wait for Clk_period;
		Addr <=  "0010010011111";
		Trees_din <= x"33058708";
		wait for Clk_period;
		Addr <=  "0010010100000";
		Trees_din <= x"0605ce04";
		wait for Clk_period;
		Addr <=  "0010010100001";
		Trees_din <= x"ff7f12e5";
		wait for Clk_period;
		Addr <=  "0010010100010";
		Trees_din <= x"fffb12e5";
		wait for Clk_period;
		Addr <=  "0010010100011";
		Trees_din <= x"9e065108";
		wait for Clk_period;
		Addr <=  "0010010100100";
		Trees_din <= x"2a063b04";
		wait for Clk_period;
		Addr <=  "0010010100101";
		Trees_din <= x"ffb012e5";
		wait for Clk_period;
		Addr <=  "0010010100110";
		Trees_din <= x"000312e5";
		wait for Clk_period;
		Addr <=  "0010010100111";
		Trees_din <= x"0302a204";
		wait for Clk_period;
		Addr <=  "0010010101000";
		Trees_din <= x"005a12e5";
		wait for Clk_period;
		Addr <=  "0010010101001";
		Trees_din <= x"fff912e5";
		wait for Clk_period;
		Addr <=  "0010010101010";
		Trees_din <= x"5200bc14";
		wait for Clk_period;
		Addr <=  "0010010101011";
		Trees_din <= x"cd010f04";
		wait for Clk_period;
		Addr <=  "0010010101100";
		Trees_din <= x"ffe712e5";
		wait for Clk_period;
		Addr <=  "0010010101101";
		Trees_din <= x"3703280c";
		wait for Clk_period;
		Addr <=  "0010010101110";
		Trees_din <= x"e5035c08";
		wait for Clk_period;
		Addr <=  "0010010101111";
		Trees_din <= x"f500ac04";
		wait for Clk_period;
		Addr <=  "0010010110000";
		Trees_din <= x"002512e5";
		wait for Clk_period;
		Addr <=  "0010010110001";
		Trees_din <= x"008912e5";
		wait for Clk_period;
		Addr <=  "0010010110010";
		Trees_din <= x"001912e5";
		wait for Clk_period;
		Addr <=  "0010010110011";
		Trees_din <= x"000b12e5";
		wait for Clk_period;
		Addr <=  "0010010110100";
		Trees_din <= x"0e03ff04";
		wait for Clk_period;
		Addr <=  "0010010110101";
		Trees_din <= x"ff9912e5";
		wait for Clk_period;
		Addr <=  "0010010110110";
		Trees_din <= x"c501bf04";
		wait for Clk_period;
		Addr <=  "0010010110111";
		Trees_din <= x"004b12e5";
		wait for Clk_period;
		Addr <=  "0010010111000";
		Trees_din <= x"ffe512e5";
		wait for Clk_period;
		Addr <=  "0010010111001";
		Trees_din <= x"6d042114";
		wait for Clk_period;
		Addr <=  "0010010111010";
		Trees_din <= x"63001f08";
		wait for Clk_period;
		Addr <=  "0010010111011";
		Trees_din <= x"5a009204";
		wait for Clk_period;
		Addr <=  "0010010111100";
		Trees_din <= x"004b1351";
		wait for Clk_period;
		Addr <=  "0010010111101";
		Trees_din <= x"ffda1351";
		wait for Clk_period;
		Addr <=  "0010010111110";
		Trees_din <= x"0607f008";
		wait for Clk_period;
		Addr <=  "0010010111111";
		Trees_din <= x"b4063b04";
		wait for Clk_period;
		Addr <=  "0010011000000";
		Trees_din <= x"ff7d1351";
		wait for Clk_period;
		Addr <=  "0010011000001";
		Trees_din <= x"ffdf1351";
		wait for Clk_period;
		Addr <=  "0010011000010";
		Trees_din <= x"fff91351";
		wait for Clk_period;
		Addr <=  "0010011000011";
		Trees_din <= x"0604b114";
		wait for Clk_period;
		Addr <=  "0010011000100";
		Trees_din <= x"33057308";
		wait for Clk_period;
		Addr <=  "0010011000101";
		Trees_din <= x"f2052e04";
		wait for Clk_period;
		Addr <=  "0010011000110";
		Trees_din <= x"ffa01351";
		wait for Clk_period;
		Addr <=  "0010011000111";
		Trees_din <= x"00011351";
		wait for Clk_period;
		Addr <=  "0010011001000";
		Trees_din <= x"d300ff08";
		wait for Clk_period;
		Addr <=  "0010011001001";
		Trees_din <= x"2d033204";
		wait for Clk_period;
		Addr <=  "0010011001010";
		Trees_din <= x"00561351";
		wait for Clk_period;
		Addr <=  "0010011001011";
		Trees_din <= x"00021351";
		wait for Clk_period;
		Addr <=  "0010011001100";
		Trees_din <= x"ffd61351";
		wait for Clk_period;
		Addr <=  "0010011001101";
		Trees_din <= x"07035d0c";
		wait for Clk_period;
		Addr <=  "0010011001110";
		Trees_din <= x"5100c804";
		wait for Clk_period;
		Addr <=  "0010011001111";
		Trees_din <= x"fff71351";
		wait for Clk_period;
		Addr <=  "0010011010000";
		Trees_din <= x"70033604";
		wait for Clk_period;
		Addr <=  "0010011010001";
		Trees_din <= x"00811351";
		wait for Clk_period;
		Addr <=  "0010011010010";
		Trees_din <= x"001f1351";
		wait for Clk_period;
		Addr <=  "0010011010011";
		Trees_din <= x"ffe51351";
		wait for Clk_period;
		Addr <=  "0010011010100";
		Trees_din <= x"15042318";
		wait for Clk_period;
		Addr <=  "0010011010101";
		Trees_din <= x"2a06640c";
		wait for Clk_period;
		Addr <=  "0010011010110";
		Trees_din <= x"240a7208";
		wait for Clk_period;
		Addr <=  "0010011010111";
		Trees_din <= x"c7000d04";
		wait for Clk_period;
		Addr <=  "0010011011000";
		Trees_din <= x"ffe613ad";
		wait for Clk_period;
		Addr <=  "0010011011001";
		Trees_din <= x"ff7f13ad";
		wait for Clk_period;
		Addr <=  "0010011011010";
		Trees_din <= x"fffe13ad";
		wait for Clk_period;
		Addr <=  "0010011011011";
		Trees_din <= x"68018b08";
		wait for Clk_period;
		Addr <=  "0010011011100";
		Trees_din <= x"24088404";
		wait for Clk_period;
		Addr <=  "0010011011101";
		Trees_din <= x"001313ad";
		wait for Clk_period;
		Addr <=  "0010011011110";
		Trees_din <= x"004613ad";
		wait for Clk_period;
		Addr <=  "0010011011111";
		Trees_din <= x"ffd013ad";
		wait for Clk_period;
		Addr <=  "0010011100000";
		Trees_din <= x"5901cf10";
		wait for Clk_period;
		Addr <=  "0010011100001";
		Trees_din <= x"cd010f04";
		wait for Clk_period;
		Addr <=  "0010011100010";
		Trees_din <= x"ffdc13ad";
		wait for Clk_period;
		Addr <=  "0010011100011";
		Trees_din <= x"5b038908";
		wait for Clk_period;
		Addr <=  "0010011100100";
		Trees_din <= x"5703cf04";
		wait for Clk_period;
		Addr <=  "0010011100101";
		Trees_din <= x"007a13ad";
		wait for Clk_period;
		Addr <=  "0010011100110";
		Trees_din <= x"001413ad";
		wait for Clk_period;
		Addr <=  "0010011100111";
		Trees_din <= x"fffa13ad";
		wait for Clk_period;
		Addr <=  "0010011101000";
		Trees_din <= x"0e063504";
		wait for Clk_period;
		Addr <=  "0010011101001";
		Trees_din <= x"ffa013ad";
		wait for Clk_period;
		Addr <=  "0010011101010";
		Trees_din <= x"001a13ad";
		wait for Clk_period;
		Addr <=  "0010011101011";
		Trees_din <= x"2803400c";
		wait for Clk_period;
		Addr <=  "0010011101100";
		Trees_din <= x"0605ce08";
		wait for Clk_period;
		Addr <=  "0010011101101";
		Trees_din <= x"24083504";
		wait for Clk_period;
		Addr <=  "0010011101110";
		Trees_din <= x"ff8913f9";
		wait for Clk_period;
		Addr <=  "0010011101111";
		Trees_din <= x"ffde13f9";
		wait for Clk_period;
		Addr <=  "0010011110000";
		Trees_din <= x"000413f9";
		wait for Clk_period;
		Addr <=  "0010011110001";
		Trees_din <= x"0e034f08";
		wait for Clk_period;
		Addr <=  "0010011110010";
		Trees_din <= x"e5018b04";
		wait for Clk_period;
		Addr <=  "0010011110011";
		Trees_din <= x"001513f9";
		wait for Clk_period;
		Addr <=  "0010011110100";
		Trees_din <= x"ff9f13f9";
		wait for Clk_period;
		Addr <=  "0010011110101";
		Trees_din <= x"0b057a10";
		wait for Clk_period;
		Addr <=  "0010011110110";
		Trees_din <= x"5902090c";
		wait for Clk_period;
		Addr <=  "0010011110111";
		Trees_din <= x"69008204";
		wait for Clk_period;
		Addr <=  "0010011111000";
		Trees_din <= x"000913f9";
		wait for Clk_period;
		Addr <=  "0010011111001";
		Trees_din <= x"0d045304";
		wait for Clk_period;
		Addr <=  "0010011111010";
		Trees_din <= x"007e13f9";
		wait for Clk_period;
		Addr <=  "0010011111011";
		Trees_din <= x"001813f9";
		wait for Clk_period;
		Addr <=  "0010011111100";
		Trees_din <= x"fff613f9";
		wait for Clk_period;
		Addr <=  "0010011111101";
		Trees_din <= x"ffdd13f9";
		wait for Clk_period;
		Addr <=  "0010011111110";
		Trees_din <= x"0a070218";
		wait for Clk_period;
		Addr <=  "0010011111111";
		Trees_din <= x"00016810";
		wait for Clk_period;
		Addr <=  "0010100000000";
		Trees_din <= x"df01aa08";
		wait for Clk_period;
		Addr <=  "0010100000001";
		Trees_din <= x"57028404";
		wait for Clk_period;
		Addr <=  "0010100000010";
		Trees_din <= x"0052144d";
		wait for Clk_period;
		Addr <=  "0010100000011";
		Trees_din <= x"ffdd144d";
		wait for Clk_period;
		Addr <=  "0010100000100";
		Trees_din <= x"1e06ea04";
		wait for Clk_period;
		Addr <=  "0010100000101";
		Trees_din <= x"ffa9144d";
		wait for Clk_period;
		Addr <=  "0010100000110";
		Trees_din <= x"000f144d";
		wait for Clk_period;
		Addr <=  "0010100000111";
		Trees_din <= x"3b010304";
		wait for Clk_period;
		Addr <=  "0010100001000";
		Trees_din <= x"ffe0144d";
		wait for Clk_period;
		Addr <=  "0010100001001";
		Trees_din <= x"ff8d144d";
		wait for Clk_period;
		Addr <=  "0010100001010";
		Trees_din <= x"b603650c";
		wait for Clk_period;
		Addr <=  "0010100001011";
		Trees_din <= x"3702b608";
		wait for Clk_period;
		Addr <=  "0010100001100";
		Trees_din <= x"df026b04";
		wait for Clk_period;
		Addr <=  "0010100001101";
		Trees_din <= x"0071144d";
		wait for Clk_period;
		Addr <=  "0010100001110";
		Trees_din <= x"001c144d";
		wait for Clk_period;
		Addr <=  "0010100001111";
		Trees_din <= x"fffe144d";
		wait for Clk_period;
		Addr <=  "0010100010000";
		Trees_din <= x"1d067a04";
		wait for Clk_period;
		Addr <=  "0010100010001";
		Trees_din <= x"ffbe144d";
		wait for Clk_period;
		Addr <=  "0010100010010";
		Trees_din <= x"0023144d";
		wait for Clk_period;
		Addr <=  "0010100010011";
		Trees_din <= x"2a05810c";
		wait for Clk_period;
		Addr <=  "0010100010100";
		Trees_din <= x"03004304";
		wait for Clk_period;
		Addr <=  "0010100010101";
		Trees_din <= x"001a1489";
		wait for Clk_period;
		Addr <=  "0010100010110";
		Trees_din <= x"6d08c404";
		wait for Clk_period;
		Addr <=  "0010100010111";
		Trees_din <= x"ff941489";
		wait for Clk_period;
		Addr <=  "0010100011000";
		Trees_din <= x"fffa1489";
		wait for Clk_period;
		Addr <=  "0010100011001";
		Trees_din <= x"0e05620c";
		wait for Clk_period;
		Addr <=  "0010100011010";
		Trees_din <= x"37010704";
		wait for Clk_period;
		Addr <=  "0010100011011";
		Trees_din <= x"002c1489";
		wait for Clk_period;
		Addr <=  "0010100011100";
		Trees_din <= x"23069904";
		wait for Clk_period;
		Addr <=  "0010100011101";
		Trees_din <= x"ffb01489";
		wait for Clk_period;
		Addr <=  "0010100011110";
		Trees_din <= x"000b1489";
		wait for Clk_period;
		Addr <=  "0010100011111";
		Trees_din <= x"1e048404";
		wait for Clk_period;
		Addr <=  "0010100100000";
		Trees_din <= x"fffd1489";
		wait for Clk_period;
		Addr <=  "0010100100001";
		Trees_din <= x"00681489";
		wait for Clk_period;
		Addr <=  "0010100100010";
		Trees_din <= x"0604b110";
		wait for Clk_period;
		Addr <=  "0010100100011";
		Trees_din <= x"5f088a08";
		wait for Clk_period;
		Addr <=  "0010100100100";
		Trees_din <= x"15042304";
		wait for Clk_period;
		Addr <=  "0010100100101";
		Trees_din <= x"ff9714cd";
		wait for Clk_period;
		Addr <=  "0010100100110";
		Trees_din <= x"fffd14cd";
		wait for Clk_period;
		Addr <=  "0010100100111";
		Trees_din <= x"53047604";
		wait for Clk_period;
		Addr <=  "0010100101000";
		Trees_din <= x"fff614cd";
		wait for Clk_period;
		Addr <=  "0010100101001";
		Trees_din <= x"002a14cd";
		wait for Clk_period;
		Addr <=  "0010100101010";
		Trees_din <= x"e701bf08";
		wait for Clk_period;
		Addr <=  "0010100101011";
		Trees_din <= x"5c014904";
		wait for Clk_period;
		Addr <=  "0010100101100";
		Trees_din <= x"002514cd";
		wait for Clk_period;
		Addr <=  "0010100101101";
		Trees_din <= x"ffbf14cd";
		wait for Clk_period;
		Addr <=  "0010100101110";
		Trees_din <= x"ee082708";
		wait for Clk_period;
		Addr <=  "0010100101111";
		Trees_din <= x"7002a304";
		wait for Clk_period;
		Addr <=  "0010100110000";
		Trees_din <= x"007014cd";
		wait for Clk_period;
		Addr <=  "0010100110001";
		Trees_din <= x"001a14cd";
		wait for Clk_period;
		Addr <=  "0010100110010";
		Trees_din <= x"ffed14cd";
		wait for Clk_period;
		Addr <=  "0010100110011";
		Trees_din <= x"33051710";
		wait for Clk_period;
		Addr <=  "0010100110100";
		Trees_din <= x"63001c08";
		wait for Clk_period;
		Addr <=  "0010100110101";
		Trees_din <= x"9300ff04";
		wait for Clk_period;
		Addr <=  "0010100110110";
		Trees_din <= x"fff51509";
		wait for Clk_period;
		Addr <=  "0010100110111";
		Trees_din <= x"003e1509";
		wait for Clk_period;
		Addr <=  "0010100111000";
		Trees_din <= x"9e083f04";
		wait for Clk_period;
		Addr <=  "0010100111001";
		Trees_din <= x"ffa01509";
		wait for Clk_period;
		Addr <=  "0010100111010";
		Trees_din <= x"00001509";
		wait for Clk_period;
		Addr <=  "0010100111011";
		Trees_din <= x"1e046004";
		wait for Clk_period;
		Addr <=  "0010100111100";
		Trees_din <= x"ffe31509";
		wait for Clk_period;
		Addr <=  "0010100111101";
		Trees_din <= x"3d01c508";
		wait for Clk_period;
		Addr <=  "0010100111110";
		Trees_din <= x"51010c04";
		wait for Clk_period;
		Addr <=  "0010100111111";
		Trees_din <= x"000f1509";
		wait for Clk_period;
		Addr <=  "0010101000000";
		Trees_din <= x"00601509";
		wait for Clk_period;
		Addr <=  "0010101000001";
		Trees_din <= x"fff51509";
		wait for Clk_period;
		Addr <=  "0010101000010";
		Trees_din <= x"1504230c";
		wait for Clk_period;
		Addr <=  "0010101000011";
		Trees_din <= x"240a7208";
		wait for Clk_period;
		Addr <=  "0010101000100";
		Trees_din <= x"2a06bb04";
		wait for Clk_period;
		Addr <=  "0010101000101";
		Trees_din <= x"ff9e153d";
		wait for Clk_period;
		Addr <=  "0010101000110";
		Trees_din <= x"fffb153d";
		wait for Clk_period;
		Addr <=  "0010101000111";
		Trees_din <= x"0018153d";
		wait for Clk_period;
		Addr <=  "0010101001000";
		Trees_din <= x"2f023108";
		wait for Clk_period;
		Addr <=  "0010101001001";
		Trees_din <= x"c402b804";
		wait for Clk_period;
		Addr <=  "0010101001010";
		Trees_din <= x"005d153d";
		wait for Clk_period;
		Addr <=  "0010101001011";
		Trees_din <= x"0001153d";
		wait for Clk_period;
		Addr <=  "0010101001100";
		Trees_din <= x"fe014f04";
		wait for Clk_period;
		Addr <=  "0010101001101";
		Trees_din <= x"001e153d";
		wait for Clk_period;
		Addr <=  "0010101001110";
		Trees_din <= x"ffc6153d";
		wait for Clk_period;
		Addr <=  "0010101001111";
		Trees_din <= x"0a04fa0c";
		wait for Clk_period;
		Addr <=  "0010101010000";
		Trees_din <= x"3306ac08";
		wait for Clk_period;
		Addr <=  "0010101010001";
		Trees_din <= x"f0007704";
		wait for Clk_period;
		Addr <=  "0010101010010";
		Trees_din <= x"fff61571";
		wait for Clk_period;
		Addr <=  "0010101010011";
		Trees_din <= x"ffa21571";
		wait for Clk_period;
		Addr <=  "0010101010100";
		Trees_din <= x"000c1571";
		wait for Clk_period;
		Addr <=  "0010101010101";
		Trees_din <= x"c502990c";
		wait for Clk_period;
		Addr <=  "0010101010110";
		Trees_din <= x"9104e204";
		wait for Clk_period;
		Addr <=  "0010101010111";
		Trees_din <= x"00031571";
		wait for Clk_period;
		Addr <=  "0010101011000";
		Trees_din <= x"1f031b04";
		wait for Clk_period;
		Addr <=  "0010101011001";
		Trees_din <= x"00161571";
		wait for Clk_period;
		Addr <=  "0010101011010";
		Trees_din <= x"005d1571";
		wait for Clk_period;
		Addr <=  "0010101011011";
		Trees_din <= x"ffe21571";
		wait for Clk_period;
		Addr <=  "0010101011100";
		Trees_din <= x"28034008";
		wait for Clk_period;
		Addr <=  "0010101011101";
		Trees_din <= x"0605ce04";
		wait for Clk_period;
		Addr <=  "0010101011110";
		Trees_din <= x"ffad15a5";
		wait for Clk_period;
		Addr <=  "0010101011111";
		Trees_din <= x"000115a5";
		wait for Clk_period;
		Addr <=  "0010101100000";
		Trees_din <= x"7604c40c";
		wait for Clk_period;
		Addr <=  "0010101100001";
		Trees_din <= x"0301cf08";
		wait for Clk_period;
		Addr <=  "0010101100010";
		Trees_din <= x"a8023804";
		wait for Clk_period;
		Addr <=  "0010101100011";
		Trees_din <= x"ffdc15a5";
		wait for Clk_period;
		Addr <=  "0010101100100";
		Trees_din <= x"003815a5";
		wait for Clk_period;
		Addr <=  "0010101100101";
		Trees_din <= x"ffbc15a5";
		wait for Clk_period;
		Addr <=  "0010101100110";
		Trees_din <= x"d3017c04";
		wait for Clk_period;
		Addr <=  "0010101100111";
		Trees_din <= x"005515a5";
		wait for Clk_period;
		Addr <=  "0010101101000";
		Trees_din <= x"000815a5";
		wait for Clk_period;
		Addr <=  "0010101101001";
		Trees_din <= x"0604b10c";
		wait for Clk_period;
		Addr <=  "0010101101010";
		Trees_din <= x"1e07f908";
		wait for Clk_period;
		Addr <=  "0010101101011";
		Trees_din <= x"15042304";
		wait for Clk_period;
		Addr <=  "0010101101100";
		Trees_din <= x"ffaa15d1";
		wait for Clk_period;
		Addr <=  "0010101101101";
		Trees_din <= x"fff815d1";
		wait for Clk_period;
		Addr <=  "0010101101110";
		Trees_din <= x"001415d1";
		wait for Clk_period;
		Addr <=  "0010101101111";
		Trees_din <= x"a2020a04";
		wait for Clk_period;
		Addr <=  "0010101110000";
		Trees_din <= x"ffe715d1";
		wait for Clk_period;
		Addr <=  "0010101110001";
		Trees_din <= x"72020604";
		wait for Clk_period;
		Addr <=  "0010101110010";
		Trees_din <= x"005215d1";
		wait for Clk_period;
		Addr <=  "0010101110011";
		Trees_din <= x"000315d1";
		wait for Clk_period;
		Addr <=  "0010101110100";
		Trees_din <= x"38035404";
		wait for Clk_period;
		Addr <=  "0010101110101";
		Trees_din <= x"ffb715fd";
		wait for Clk_period;
		Addr <=  "0010101110110";
		Trees_din <= x"5e02720c";
		wait for Clk_period;
		Addr <=  "0010101110111";
		Trees_din <= x"0b039508";
		wait for Clk_period;
		Addr <=  "0010101111000";
		Trees_din <= x"be004704";
		wait for Clk_period;
		Addr <=  "0010101111001";
		Trees_din <= x"000a15fd";
		wait for Clk_period;
		Addr <=  "0010101111010";
		Trees_din <= x"005915fd";
		wait for Clk_period;
		Addr <=  "0010101111011";
		Trees_din <= x"fff715fd";
		wait for Clk_period;
		Addr <=  "0010101111100";
		Trees_din <= x"c903e504";
		wait for Clk_period;
		Addr <=  "0010101111101";
		Trees_din <= x"ffc915fd";
		wait for Clk_period;
		Addr <=  "0010101111110";
		Trees_din <= x"000d15fd";
		wait for Clk_period;
		Addr <=  "0010101111111";
		Trees_din <= x"0a07020c";
		wait for Clk_period;
		Addr <=  "0010110000000";
		Trees_din <= x"3b010d04";
		wait for Clk_period;
		Addr <=  "0010110000001";
		Trees_din <= x"000b1629";
		wait for Clk_period;
		Addr <=  "0010110000010";
		Trees_din <= x"f000b404";
		wait for Clk_period;
		Addr <=  "0010110000011";
		Trees_din <= x"fff41629";
		wait for Clk_period;
		Addr <=  "0010110000100";
		Trees_din <= x"ffaf1629";
		wait for Clk_period;
		Addr <=  "0010110000101";
		Trees_din <= x"3504e708";
		wait for Clk_period;
		Addr <=  "0010110000110";
		Trees_din <= x"2e010d04";
		wait for Clk_period;
		Addr <=  "0010110000111";
		Trees_din <= x"00511629";
		wait for Clk_period;
		Addr <=  "0010110001000";
		Trees_din <= x"00091629";
		wait for Clk_period;
		Addr <=  "0010110001001";
		Trees_din <= x"fff01629";
		wait for Clk_period;
		Addr <=  "0010110001010";
		Trees_din <= x"28034008";
		wait for Clk_period;
		Addr <=  "0010110001011";
		Trees_din <= x"d6021d04";
		wait for Clk_period;
		Addr <=  "0010110001100";
		Trees_din <= x"fff2165d";
		wait for Clk_period;
		Addr <=  "0010110001101";
		Trees_din <= x"ffb6165d";
		wait for Clk_period;
		Addr <=  "0010110001110";
		Trees_din <= x"1802d70c";
		wait for Clk_period;
		Addr <=  "0010110001111";
		Trees_din <= x"e0006d04";
		wait for Clk_period;
		Addr <=  "0010110010000";
		Trees_din <= x"0002165d";
		wait for Clk_period;
		Addr <=  "0010110010001";
		Trees_din <= x"1503da04";
		wait for Clk_period;
		Addr <=  "0010110010010";
		Trees_din <= x"0015165d";
		wait for Clk_period;
		Addr <=  "0010110010011";
		Trees_din <= x"0058165d";
		wait for Clk_period;
		Addr <=  "0010110010100";
		Trees_din <= x"0301cf04";
		wait for Clk_period;
		Addr <=  "0010110010101";
		Trees_din <= x"000e165d";
		wait for Clk_period;
		Addr <=  "0010110010110";
		Trees_din <= x"ffc9165d";
		wait for Clk_period;
		Addr <=  "0010110010111";
		Trees_din <= x"df02020c";
		wait for Clk_period;
		Addr <=  "0010110011000";
		Trees_din <= x"3702f908";
		wait for Clk_period;
		Addr <=  "0010110011001";
		Trees_din <= x"5e024104";
		wait for Clk_period;
		Addr <=  "0010110011010";
		Trees_din <= x"004d1681";
		wait for Clk_period;
		Addr <=  "0010110011011";
		Trees_din <= x"00041681";
		wait for Clk_period;
		Addr <=  "0010110011100";
		Trees_din <= x"ffdd1681";
		wait for Clk_period;
		Addr <=  "0010110011101";
		Trees_din <= x"2407ce04";
		wait for Clk_period;
		Addr <=  "0010110011110";
		Trees_din <= x"ffbe1681";
		wait for Clk_period;
		Addr <=  "0010110011111";
		Trees_din <= x"00081681";
		wait for Clk_period;
		Addr <=  "0010110100000";
		Trees_din <= x"0604b10c";
		wait for Clk_period;
		Addr <=  "0010110100001";
		Trees_din <= x"73067008";
		wait for Clk_period;
		Addr <=  "0010110100010";
		Trees_din <= x"9d00ef04";
		wait for Clk_period;
		Addr <=  "0010110100011";
		Trees_din <= x"fff216ad";
		wait for Clk_period;
		Addr <=  "0010110100100";
		Trees_din <= x"ffb416ad";
		wait for Clk_period;
		Addr <=  "0010110100101";
		Trees_din <= x"000c16ad";
		wait for Clk_period;
		Addr <=  "0010110100110";
		Trees_din <= x"a2020a04";
		wait for Clk_period;
		Addr <=  "0010110100111";
		Trees_din <= x"ffec16ad";
		wait for Clk_period;
		Addr <=  "0010110101000";
		Trees_din <= x"35040404";
		wait for Clk_period;
		Addr <=  "0010110101001";
		Trees_din <= x"004716ad";
		wait for Clk_period;
		Addr <=  "0010110101010";
		Trees_din <= x"000d16ad";
		wait for Clk_period;
		Addr <=  "0010110101011";
		Trees_din <= x"3305320c";
		wait for Clk_period;
		Addr <=  "0010110101100";
		Trees_din <= x"63001c04";
		wait for Clk_period;
		Addr <=  "0010110101101";
		Trees_din <= x"001316d9";
		wait for Clk_period;
		Addr <=  "0010110101110";
		Trees_din <= x"4e062004";
		wait for Clk_period;
		Addr <=  "0010110101111";
		Trees_din <= x"ffb916d9";
		wait for Clk_period;
		Addr <=  "0010110110000";
		Trees_din <= x"ffee16d9";
		wait for Clk_period;
		Addr <=  "0010110110001";
		Trees_din <= x"70029b08";
		wait for Clk_period;
		Addr <=  "0010110110010";
		Trees_din <= x"28050e04";
		wait for Clk_period;
		Addr <=  "0010110110011";
		Trees_din <= x"000516d9";
		wait for Clk_period;
		Addr <=  "0010110110100";
		Trees_din <= x"004916d9";
		wait for Clk_period;
		Addr <=  "0010110110101";
		Trees_din <= x"fff116d9";
		wait for Clk_period;
		Addr <=  "0010110110110";
		Trees_din <= x"2a058108";
		wait for Clk_period;
		Addr <=  "0010110110111";
		Trees_din <= x"0b023704";
		wait for Clk_period;
		Addr <=  "0010110111000";
		Trees_din <= x"000916fd";
		wait for Clk_period;
		Addr <=  "0010110111001";
		Trees_din <= x"ffbf16fd";
		wait for Clk_period;
		Addr <=  "0010110111010";
		Trees_din <= x"72020608";
		wait for Clk_period;
		Addr <=  "0010110111011";
		Trees_din <= x"a2020504";
		wait for Clk_period;
		Addr <=  "0010110111100";
		Trees_din <= x"fffe16fd";
		wait for Clk_period;
		Addr <=  "0010110111101";
		Trees_din <= x"004716fd";
		wait for Clk_period;
		Addr <=  "0010110111110";
		Trees_din <= x"ffe616fd";
		wait for Clk_period;
		Addr <=  "0010110111111";
		Trees_din <= x"06034708";
		wait for Clk_period;
		Addr <=  "0010111000000";
		Trees_din <= x"9d010804";
		wait for Clk_period;
		Addr <=  "0010111000001";
		Trees_din <= x"fff61729";
		wait for Clk_period;
		Addr <=  "0010111000010";
		Trees_din <= x"ffc81729";
		wait for Clk_period;
		Addr <=  "0010111000011";
		Trees_din <= x"1f048308";
		wait for Clk_period;
		Addr <=  "0010111000100";
		Trees_din <= x"37016f04";
		wait for Clk_period;
		Addr <=  "0010111000101";
		Trees_din <= x"00191729";
		wait for Clk_period;
		Addr <=  "0010111000110";
		Trees_din <= x"ffd71729";
		wait for Clk_period;
		Addr <=  "0010111000111";
		Trees_din <= x"2a065604";
		wait for Clk_period;
		Addr <=  "0010111001000";
		Trees_din <= x"00101729";
		wait for Clk_period;
		Addr <=  "0010111001001";
		Trees_din <= x"00421729";
		wait for Clk_period;
		Addr <=  "0010111001010";
		Trees_din <= x"2804d108";
		wait for Clk_period;
		Addr <=  "0010111001011";
		Trees_din <= x"0000a804";
		wait for Clk_period;
		Addr <=  "0010111001100";
		Trees_din <= x"00091745";
		wait for Clk_period;
		Addr <=  "0010111001101";
		Trees_din <= x"ffc41745";
		wait for Clk_period;
		Addr <=  "0010111001110";
		Trees_din <= x"1802d704";
		wait for Clk_period;
		Addr <=  "0010111001111";
		Trees_din <= x"00371745";
		wait for Clk_period;
		Addr <=  "0010111010000";
		Trees_din <= x"fff31745";
		wait for Clk_period;
		Addr <=  "0010111010001";
		Trees_din <= x"0a02d804";
		wait for Clk_period;
		Addr <=  "0010111010010";
		Trees_din <= x"ffcd1761";
		wait for Clk_period;
		Addr <=  "0010111010011";
		Trees_din <= x"1f03b804";
		wait for Clk_period;
		Addr <=  "0010111010100";
		Trees_din <= x"ffec1761";
		wait for Clk_period;
		Addr <=  "0010111010101";
		Trees_din <= x"9105d404";
		wait for Clk_period;
		Addr <=  "0010111010110";
		Trees_din <= x"00011761";
		wait for Clk_period;
		Addr <=  "0010111010111";
		Trees_din <= x"00421761";
		wait for Clk_period;
		Addr <=  "0010111011000";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  1
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"51015b38";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"23072524";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"4a00f414";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"c001410c";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"37007b04";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"ff8900f5";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"6900a204";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"039200f5";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"008e00f5";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"07045604";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"ff6400f5";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"013c00f5";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"c004b80c";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"8703db08";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"cb00f904";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"ff9d00f5";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"042b00f5";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"000000f5";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"ffe500f5";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"8701710c";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"cb032908";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"2f02a404";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"ff7d00f5";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"01c600f5";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"037900f5";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"99000b04";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"01c600f5";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"ff5900f5";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"a601231c";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"6f007b08";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"0c02e104";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"ff6700f5";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"00b200f5";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"f7012f08";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"02037b04";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"00b200f5";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"ff8900f5";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"14003204";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"001200f5";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"67061004";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"03f400f5";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"013c00f5";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"6500260c";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"cc00e808";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"0102ec04";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"ff8900f5";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"002700f5";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"033200f5";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"6900990c";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"99003804";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"02dc00f5";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"8700d004";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"015400f5";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"ff7200f5";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"93000a08";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"07033a04";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"ff7300f5";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"01c600f5";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"ec001204";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"002700f5";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"ff4e00f5";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"5101ef3c";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"7607ed30";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"2c007710";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"b3021b08";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"26018a04";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"ff5501c1";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"003201c1";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"69007204";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"017101c1";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"ff9001c1";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"0c006a10";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"bb00fa08";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"93006904";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"019301c1";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"ffa901c1";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"f4002404";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"00ab01c1";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"ff5901c1";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"d5019c08";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"050d8704";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"01a901c1";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"ff8101c1";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"77040704";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"ff6e01c1";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"00b101c1";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"ef016c04";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"ff5901c1";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"a6020c04";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"012301c1";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"ff8601c1";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"a6014714";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"65015510";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"2c011604";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"ff8701c1";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"3b009b04";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"ff9e01c1";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"3000cf04";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"000701c1";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"01a301c1";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"ff6c01c1";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"c8004708";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"5c023304";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"ff7b01c1";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"015801c1";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"2500e70c";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"2902f304";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"ff6c01c1";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"08025204";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"003901c1";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"014a01c1";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"ff5401c1";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"5101ef44";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"87024928";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"c004b820";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"0c004410";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"6f016708";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"93000604";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"007f029d";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"ff55029d";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"d5007e04";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"012f029d";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"ff95029d";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"4a008608";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"f3038004";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"ff6b029d";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"00c0029d";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"37003d04";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"008d029d";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"0131029d";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"9809dd04";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"ff69029d";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"003b029d";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"26020110";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"1404aa08";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"5a070004";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"ff59029d";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"0018029d";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"43014804";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"ff99029d";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"0136029d";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"d500a608";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"3a020d04";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"0003029d";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"012f029d";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"ff7d029d";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"99003118";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"8600ec08";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"71010304";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"0022029d";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"ff67029d";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"6f006204";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"ff86029d";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"0c006a04";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"ff90029d";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"9c00cc04";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"0038029d";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"0146029d";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"a600a108";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"40007304";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"00c0029d";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"0023029d";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"65001e04";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"0028029d";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"81001b04";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"fff7029d";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"ff58029d";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"69014234";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"c0042124";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"0e056214";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"2c003b08";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"7a016204";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"ff720359";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"00220359";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"93038e08";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"3000cf04";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"007d0359";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"00f80359";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"ff790359";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"2601d808";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"cd010804";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"00920359";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"ff540359";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"be005704";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"00fc0359";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"ff870359";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"49048b08";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"48039504";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"ff620359";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"000d0359";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"12007904";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"00cd0359";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"00080359";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"51011810";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"ef00a004";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"ff5f0359";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"ca017508";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"a7022404";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"00060359";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"00f90359";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"ff8f0359";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"2500ea0c";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"6201d104";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"ff7d0359";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"7f00ec04";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"001a0359";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"00f30359";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"8a08210c";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"be000004";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"00340359";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"fc000004";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"00160359";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"ff5b0359";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"00820359";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"6501364c";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"5200441c";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"6900da14";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"29012508";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"7403c604";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"ff5a041d";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"0080041d";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"b601b908";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"da002904";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"ff66041d";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"0088041d";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"00dd041d";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"ad051704";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"ff5e041d";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"0006041d";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"fc03e71c";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"6e00760c";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"77012d04";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"ff3b041d";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"37009604";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"ffa3041d";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"00c7041d";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"a80a3808";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"ac080d04";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"00d8041d";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"ff94041d";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"0903a004";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"ff70041d";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"0090041d";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"c4027d08";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"33025c04";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"006b041d";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"ff62041d";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"c0014108";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"1a00fd04";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"0027041d";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"00d0041d";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"ffa8041d";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"2500f510";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"b1018e08";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"af015c04";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"fff5041d";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"00c9041d";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"9004bf04";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"ff71041d";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"0027041d";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"ec002804";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"000e041d";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"ff5d041d";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"6501365c";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"0c010d30";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"e600f11c";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"6200d910";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"c7010708";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"e902ec04";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"ff680501";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"ffeb0501";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"65003504";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"00a40501";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"ffe80501";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"5c005d04";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"ff860501";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"d500bb04";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"00bd0501";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"ffc00501";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"2f02f908";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"22000304";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"fff90501";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"ff460501";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"51013308";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"5400a804";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"00a20501";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"00250501";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"ff8a0501";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"24097e1c";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"2c005e0c";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"92046808";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"b9004304";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"fff70501";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"ff750501";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"00820501";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"23084c08";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"08002804";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"00350501";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"00c50501";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"6100fc04";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"007b0501";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"ff6d0501";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"b8036608";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"47031104";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"ff6c0501";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"00090501";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"6f00d104";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"ffe40501";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"00a80501";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"2500f510";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"b1018e08";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"af015c04";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"fff20501";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"00b00501";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"41025404";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"ff790501";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"00200501";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"ec002804";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"00080501";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"ff600501";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"5101ef50";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"0c015c34";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"3d016520";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"69009910";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"63002208";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"cb042f04";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"ff4c05e5";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"007905e5";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"b300ce04";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"ffae05e5";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"00b305e5";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"07021b08";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"94000e04";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"000405e5";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"ff4d05e5";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"87018f04";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"007205e5";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"ff9c05e5";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"3e05fc10";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"fe007608";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"29020804";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"ff9005e5";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"006505e5";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"9401db04";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"00bd05e5";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"002f05e5";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"ff8205e5";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"61066714";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"a603fd0c";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"2d083a08";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"07007704";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"004705e5";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"00b805e5";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"ff7b05e5";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"6e028804";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"ff7e05e5";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"006605e5";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"3b068d04";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"ffdb05e5";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"ff4c05e5";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"99003114";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"6200e704";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"ff7a05e5";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"0207f60c";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"cc010304";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"ffae05e5";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"9c00d204";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"001d05e5";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"00b605e5";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"ff8b05e5";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"a600a104";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"005c05e5";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"81001b04";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"000b05e5";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"25003804";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"fff605e5";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"ff6205e5";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"25028f54";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"4a01632c";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"6900a614";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"c001f30c";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"790b7e08";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"0c006a04";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"ffdd06c9";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"00a806c9";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"ff5706c9";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"f2031004";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"ff7506c9";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"005706c9";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"1405b010";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"6f022808";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"7704d104";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"ff6306c9";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"001306c9";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"c8011004";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"007206c9";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"ffa206c9";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"ec019e04";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"009f06c9";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"002206c9";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"d2062820";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"37003d10";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"d2015308";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"4801d404";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"008f06c9";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"002506c9";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"97022a04";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"ffdd06c9";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"ff0206c9";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"e5002308";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"5200a604";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"ff8406c9";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"004706c9";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"08002804";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"002906c9";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"00ae06c9";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"8603bf04";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"ff7606c9";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"004706c9";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"6900e614";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"e601150c";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"49016f04";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"ffc406c9";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"37010f04";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"000506c9";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"009d06c9";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"cb017d04";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"000606c9";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"ff7706c9";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"a600b004";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"003b06c9";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"ed000404";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"ffff06c9";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"ff6106c9";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"6501365c";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"26016438";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"0c01b61c";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"fa01d40c";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"b002fe04";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"ff3c07a5";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"07019304";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"ff8907a5";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"005007a5";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"9300ff08";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"ec023804";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"007207a5";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"ffb207a5";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"cd00c004";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"001607a5";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"ff4507a5";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"68024510";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"8f022a08";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"51021304";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"007807a5";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"ff9f07a5";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"b2031d04";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"ff4c07a5";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"ffce07a5";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"a4006004";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"ffb107a5";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"e0018c04";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"00a707a5";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"ffee07a5";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"6105e51c";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"23084c10";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"6e006608";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"41032404";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"ff6707a5";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"007e07a5";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"d3000904";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"ffce07a5";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"00a807a5";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"87016004";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"008107a5";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"a8023804";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"ff8207a5";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"ffdd07a5";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"0a019404";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"ff4907a5";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"006607a5";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"2500f50c";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"7400e404";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"ff9207a5";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"3a016d04";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"ffce07a5";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"008b07a5";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"ec002804";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"fff907a5";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"ff6407a5";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"25028f4c";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"2601642c";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"0c020b18";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"65000b08";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"9001a104";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"0025087d";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"0087087d";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"54007508";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"8f022a04";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"0064087d";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"ffa4087d";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"5b02fc04";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"ff3e087d";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"ffdc087d";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"8f02690c";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"51022b08";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"22009304";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"002f087d";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"00a4087d";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"ffcc087d";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"99002a04";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"0035087d";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"ff58087d";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"6105e518";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"e1043c10";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"08002808";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"3001dd04";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"ff70087d";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"007c087d";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"37002b04";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"0012087d";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"00a4087d";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"f7035c04";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"ff8c087d";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"004c087d";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"41033b04";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"ff59087d";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"005b087d";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"6900e610";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"e6011508";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"82015504";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"ffdb087d";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"007f087d";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"0002aa04";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"ff8a087d";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"fff0087d";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"a600b004";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"0028087d";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"a3071904";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"ff64087d";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"4b030b04";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"ffaf087d";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"fff0087d";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"25022354";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"4a01632c";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"0c020b18";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"1402d30c";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"65000d04";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"004d0969";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"54003304";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"00160969";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"ff690969";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"fc030a08";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"9202db04";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"00110969";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"008a0969";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"ffb70969";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"ca00be0c";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"f806a408";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"f901a904";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"00290969";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"009c0969";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"ffe50969";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"bb008304";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"00120969";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"ffa60969";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"22004910";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"2f02f008";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"58014a04";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"00080969";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"ff4b0969";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"d202d604";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"00850969";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"ffd00969";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"3b00b00c";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"c7012e04";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"ff780969";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"0c014704";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"ffd60969";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"00870969";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"f3001904";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"ffa00969";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"da026b04";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"00a10969";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"fffc0969";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"8100e318";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"6f017a10";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"8401cf08";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"a6012904";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"006a0969";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"ffc50969";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"df024904";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"ff780969";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"ffe40969";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"c001ba04";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"008e0969";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"ffdf0969";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"93008108";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"86020e04";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"ffb20969";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"00470969";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"ff630969";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"2502233c";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"3d008c1c";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"2901bb0c";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"6803b308";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"f2060a04";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"ff500a1d";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"ffe00a1d";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"000c0a1d";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"6b05570c";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"d500bb08";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"0c00c904";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"00260a1d";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"00940a1d";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"ffdb0a1d";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"ff7b0a1d";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"ec03ff18";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"6105e510";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"8a00b908";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"c601ff04";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"004b0a1d";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"ff790a1d";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"22004304";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"00190a1d";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"009c0a1d";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"17005f04";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"ff680a1d";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"003d0a1d";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"af01e404";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"ff970a1d";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"00030a1d";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"8100e314";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"f302820c";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"ef026b08";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"6403d804";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"ff800a1d";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"001c0a1d";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"005a0a1d";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"88025c04";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"000e0a1d";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"00860a1d";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"e0003204";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"fffd0a1d";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"93006904";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"ffd90a1d";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"ff620a1d";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"25020540";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"26018a28";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"7001ec14";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"fa023508";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"b0036504";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"ff4d0ad9";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"00190ad9";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"87013608";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"b1018e04";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"00810ad9";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"ffe30ad9";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"ff950ad9";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"eb01af0c";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"22002904";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"ffab0ad9";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"3b00cd04";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"fffd0ad9";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"00920ad9";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"69005b04";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"001c0ad9";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"ff970ad9";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"6105e514";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"07007708";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"c7015904";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"ff840ad9";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"005e0ad9";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"e1042b08";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"5401f604";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"009d0ad9";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"00080ad9";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"ffd80ad9";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"ffb10ad9";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"6900e614";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"2903660c";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"a7038808";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"6a00d904";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"00020ad9";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"ff620ad9";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"004c0ad9";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"93011b04";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"00840ad9";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"000f0ad9";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"a600cb04";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"002b0ad9";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"a3071904";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"ff680ad9";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"ffd30ad9";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"25020540";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"26018a24";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"0c020b14";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"fc007104";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"005b0b8d";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"99000b08";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"cf02a804";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"ffec0b8d";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"00560b8d";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"5b02b204";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"ff580b8d";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"ffd70b8d";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"8f026908";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"6b061204";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"00930b8d";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"fff40b8d";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"99002a04";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"002d0b8d";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"ff830b8d";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"da026b14";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"07007708";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"8002e404";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"ff8c0b8d";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"00530b8d";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"e1042b08";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"08002804";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"00010b8d";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"009b0b8d";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"ffdc0b8d";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"3a019d04";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"ff790b8d";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"004b0b8d";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"81010c14";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"a3021508";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"ae030e04";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"00220b8d";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"ff890b8d";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"6e012f04";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"ffe00b8d";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"f7021204";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"00210b8d";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"007f0b8d";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"93008104";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"00080b8d";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"ff670b8d";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"2501f238";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"3d008c18";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"2902e010";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"67013c08";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"13024104";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"ff350c31";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"ffdc0c31";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"4d049204";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"00400c31";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"ffb70c31";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"87013604";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"00750c31";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"fffe0c31";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"7000980c";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"66023308";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"a0002c04";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"000b0c31";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"ff830c31";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"005e0c31";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"6105e510";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"22004908";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"1f067904";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"00510c31";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"ff970c31";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"2408d604";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"00990c31";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"fff60c31";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"ffc10c31";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"f4010214";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"6f01810c";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"2902e008";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"9e022804";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"ffe20c31";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"ff850c31";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"00230c31";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"c001dc04";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"00750c31";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"ffe20c31";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"93006404";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"ffef0c31";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"ff6a0c31";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"2601642c";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"93006d14";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"fa01e208";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"5900dd04";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"ff740ce5";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"00220ce5";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"a6025e08";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"c7008004";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"00200ce5";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"00880ce5";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"ffed0ce5";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"81008a0c";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"8f016808";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"0c018b04";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"fff60ce5";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"005d0ce5";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"ffbc0ce5";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"cd012808";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"b3023c04";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"ff910ce5";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"00340ce5";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"ff690ce5";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"8701ab1c";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"da021d14";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"08002804";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"ffef0ce5";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"4a011f08";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"8700f204";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"005c0ce5";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"ffc20ce5";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"76067e04";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"009a0ce5";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"002d0ce5";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"19023e04";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"ff8e0ce5";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"003f0ce5";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"d500910c";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"e0009908";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"c4013e04";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"00220ce5";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"00790ce5";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"ffcc0ce5";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"bf009f04";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"00000ce5";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"ff880ce5";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"26016428";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"54009014";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"4100f808";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"d301f504";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"ff8f0d81";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"00030d81";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"8701ab08";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"3f01e004";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"00150d81";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"00840d81";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"ffec0d81";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"99000b08";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"f7042204";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"00530d81";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"ffe30d81";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"e7005604";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"fffe0d81";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"65001e04";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"ffe70d81";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"ff660d81";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"8701ab18";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"da021d10";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"30016b08";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"6e016404";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"ffb40d81";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"005c0d81";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"e702b004";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"00980d81";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"000e0d81";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"d200d104";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"ff980d81";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"003a0d81";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"be006408";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"5900c404";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"ffc00d81";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"006e0d81";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"b604fa04";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"ff9b0d81";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"000a0d81";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"26016b24";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"bb00ed18";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"81010c0c";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"6500bf08";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"ce01c404";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"000a0e1d";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"00780e1d";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"ffd90e1d";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"b3026704";
		wait for Clk_period;
		Addr <=  "0001101101001";
		Trees_din <= x"ff860e1d";
		wait for Clk_period;
		Addr <=  "0001101101010";
		Trees_din <= x"88023104";
		wait for Clk_period;
		Addr <=  "0001101101011";
		Trees_din <= x"ffcc0e1d";
		wait for Clk_period;
		Addr <=  "0001101101100";
		Trees_din <= x"00490e1d";
		wait for Clk_period;
		Addr <=  "0001101101101";
		Trees_din <= x"ea004d04";
		wait for Clk_period;
		Addr <=  "0001101101110";
		Trees_din <= x"fff70e1d";
		wait for Clk_period;
		Addr <=  "0001101101111";
		Trees_din <= x"a0000c04";
		wait for Clk_period;
		Addr <=  "0001101110000";
		Trees_din <= x"ffe30e1d";
		wait for Clk_period;
		Addr <=  "0001101110001";
		Trees_din <= x"ff6a0e1d";
		wait for Clk_period;
		Addr <=  "0001101110010";
		Trees_din <= x"87012d14";
		wait for Clk_period;
		Addr <=  "0001101110011";
		Trees_din <= x"da021d0c";
		wait for Clk_period;
		Addr <=  "0001101110100";
		Trees_din <= x"08002804";
		wait for Clk_period;
		Addr <=  "0001101110101";
		Trees_din <= x"ffeb0e1d";
		wait for Clk_period;
		Addr <=  "0001101110110";
		Trees_din <= x"30011504";
		wait for Clk_period;
		Addr <=  "0001101110111";
		Trees_din <= x"00250e1d";
		wait for Clk_period;
		Addr <=  "0001101111000";
		Trees_din <= x"00990e1d";
		wait for Clk_period;
		Addr <=  "0001101111001";
		Trees_din <= x"d200af04";
		wait for Clk_period;
		Addr <=  "0001101111010";
		Trees_din <= x"ffa50e1d";
		wait for Clk_period;
		Addr <=  "0001101111011";
		Trees_din <= x"002f0e1d";
		wait for Clk_period;
		Addr <=  "0001101111100";
		Trees_din <= x"94017110";
		wait for Clk_period;
		Addr <=  "0001101111101";
		Trees_din <= x"2307820c";
		wait for Clk_period;
		Addr <=  "0001101111110";
		Trees_din <= x"0e05c208";
		wait for Clk_period;
		Addr <=  "0001101111111";
		Trees_din <= x"3d00a504";
		wait for Clk_period;
		Addr <=  "0001110000000";
		Trees_din <= x"00240e1d";
		wait for Clk_period;
		Addr <=  "0001110000001";
		Trees_din <= x"007f0e1d";
		wait for Clk_period;
		Addr <=  "0001110000010";
		Trees_din <= x"fffd0e1d";
		wait for Clk_period;
		Addr <=  "0001110000011";
		Trees_din <= x"ffc40e1d";
		wait for Clk_period;
		Addr <=  "0001110000100";
		Trees_din <= x"ec015f04";
		wait for Clk_period;
		Addr <=  "0001110000101";
		Trees_din <= x"fff40e1d";
		wait for Clk_period;
		Addr <=  "0001110000110";
		Trees_din <= x"ff940e1d";
		wait for Clk_period;
		Addr <=  "0001110000111";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0001110001000";
		Trees_din <= x"26018a28";
		wait for Clk_period;
		Addr <=  "0001110001001";
		Trees_din <= x"99003a18";
		wait for Clk_period;
		Addr <=  "0001110001010";
		Trees_din <= x"0c020b10";
		wait for Clk_period;
		Addr <=  "0001110001011";
		Trees_din <= x"8e028708";
		wait for Clk_period;
		Addr <=  "0001110001100";
		Trees_din <= x"cb029f04";
		wait for Clk_period;
		Addr <=  "0001110001101";
		Trees_din <= x"ffc90ebd";
		wait for Clk_period;
		Addr <=  "0001110001110";
		Trees_din <= x"003e0ebd";
		wait for Clk_period;
		Addr <=  "0001110001111";
		Trees_din <= x"c701f804";
		wait for Clk_period;
		Addr <=  "0001110010000";
		Trees_din <= x"ffdd0ebd";
		wait for Clk_period;
		Addr <=  "0001110010001";
		Trees_din <= x"ff6c0ebd";
		wait for Clk_period;
		Addr <=  "0001110010010";
		Trees_din <= x"c0012904";
		wait for Clk_period;
		Addr <=  "0001110010011";
		Trees_din <= x"00780ebd";
		wait for Clk_period;
		Addr <=  "0001110010100";
		Trees_din <= x"00160ebd";
		wait for Clk_period;
		Addr <=  "0001110010101";
		Trees_din <= x"81007d08";
		wait for Clk_period;
		Addr <=  "0001110010110";
		Trees_din <= x"5400bd04";
		wait for Clk_period;
		Addr <=  "0001110010111";
		Trees_din <= x"003b0ebd";
		wait for Clk_period;
		Addr <=  "0001110011000";
		Trees_din <= x"ffc30ebd";
		wait for Clk_period;
		Addr <=  "0001110011001";
		Trees_din <= x"be003b04";
		wait for Clk_period;
		Addr <=  "0001110011010";
		Trees_din <= x"ffd80ebd";
		wait for Clk_period;
		Addr <=  "0001110011011";
		Trees_din <= x"ff740ebd";
		wait for Clk_period;
		Addr <=  "0001110011100";
		Trees_din <= x"da026b20";
		wait for Clk_period;
		Addr <=  "0001110011101";
		Trees_din <= x"0701030c";
		wait for Clk_period;
		Addr <=  "0001110011110";
		Trees_din <= x"9601fb04";
		wait for Clk_period;
		Addr <=  "0001110011111";
		Trees_din <= x"ffaf0ebd";
		wait for Clk_period;
		Addr <=  "0001110100000";
		Trees_din <= x"5100e804";
		wait for Clk_period;
		Addr <=  "0001110100001";
		Trees_din <= x"005f0ebd";
		wait for Clk_period;
		Addr <=  "0001110100010";
		Trees_din <= x"00080ebd";
		wait for Clk_period;
		Addr <=  "0001110100011";
		Trees_din <= x"76060c0c";
		wait for Clk_period;
		Addr <=  "0001110100100";
		Trees_din <= x"6900e604";
		wait for Clk_period;
		Addr <=  "0001110100101";
		Trees_din <= x"00970ebd";
		wait for Clk_period;
		Addr <=  "0001110100110";
		Trees_din <= x"ef029704";
		wait for Clk_period;
		Addr <=  "0001110100111";
		Trees_din <= x"00060ebd";
		wait for Clk_period;
		Addr <=  "0001110101000";
		Trees_din <= x"00530ebd";
		wait for Clk_period;
		Addr <=  "0001110101001";
		Trees_din <= x"bf009004";
		wait for Clk_period;
		Addr <=  "0001110101010";
		Trees_din <= x"003e0ebd";
		wait for Clk_period;
		Addr <=  "0001110101011";
		Trees_din <= x"ffd30ebd";
		wait for Clk_period;
		Addr <=  "0001110101100";
		Trees_din <= x"3a01b604";
		wait for Clk_period;
		Addr <=  "0001110101101";
		Trees_din <= x"ffa30ebd";
		wait for Clk_period;
		Addr <=  "0001110101110";
		Trees_din <= x"00090ebd";
		wait for Clk_period;
		Addr <=  "0001110101111";
		Trees_din <= x"26018a24";
		wait for Clk_period;
		Addr <=  "0001110110000";
		Trees_din <= x"54009010";
		wait for Clk_period;
		Addr <=  "0001110110001";
		Trees_din <= x"4100f808";
		wait for Clk_period;
		Addr <=  "0001110110010";
		Trees_din <= x"6101a004";
		wait for Clk_period;
		Addr <=  "0001110110011";
		Trees_din <= x"fff80f39";
		wait for Clk_period;
		Addr <=  "0001110110100";
		Trees_din <= x"ffa90f39";
		wait for Clk_period;
		Addr <=  "0001110110101";
		Trees_din <= x"2501e104";
		wait for Clk_period;
		Addr <=  "0001110110110";
		Trees_din <= x"006e0f39";
		wait for Clk_period;
		Addr <=  "0001110110111";
		Trees_din <= x"fffd0f39";
		wait for Clk_period;
		Addr <=  "0001110111000";
		Trees_din <= x"99000b08";
		wait for Clk_period;
		Addr <=  "0001110111001";
		Trees_din <= x"cd015a04";
		wait for Clk_period;
		Addr <=  "0001110111010";
		Trees_din <= x"00440f39";
		wait for Clk_period;
		Addr <=  "0001110111011";
		Trees_din <= x"fff40f39";
		wait for Clk_period;
		Addr <=  "0001110111100";
		Trees_din <= x"25009e04";
		wait for Clk_period;
		Addr <=  "0001110111101";
		Trees_din <= x"ffff0f39";
		wait for Clk_period;
		Addr <=  "0001110111110";
		Trees_din <= x"e7005004";
		wait for Clk_period;
		Addr <=  "0001110111111";
		Trees_din <= x"ffe70f39";
		wait for Clk_period;
		Addr <=  "0001111000000";
		Trees_din <= x"ff770f39";
		wait for Clk_period;
		Addr <=  "0001111000001";
		Trees_din <= x"2f019208";
		wait for Clk_period;
		Addr <=  "0001111000010";
		Trees_din <= x"0b03ab04";
		wait for Clk_period;
		Addr <=  "0001111000011";
		Trees_din <= x"00330f39";
		wait for Clk_period;
		Addr <=  "0001111000100";
		Trees_din <= x"ffa70f39";
		wait for Clk_period;
		Addr <=  "0001111000101";
		Trees_din <= x"87019e08";
		wait for Clk_period;
		Addr <=  "0001111000110";
		Trees_din <= x"bb01a604";
		wait for Clk_period;
		Addr <=  "0001111000111";
		Trees_din <= x"00940f39";
		wait for Clk_period;
		Addr <=  "0001111001000";
		Trees_din <= x"000f0f39";
		wait for Clk_period;
		Addr <=  "0001111001001";
		Trees_din <= x"41021504";
		wait for Clk_period;
		Addr <=  "0001111001010";
		Trees_din <= x"ffbb0f39";
		wait for Clk_period;
		Addr <=  "0001111001011";
		Trees_din <= x"bd029e04";
		wait for Clk_period;
		Addr <=  "0001111001100";
		Trees_din <= x"00050f39";
		wait for Clk_period;
		Addr <=  "0001111001101";
		Trees_din <= x"00590f39";
		wait for Clk_period;
		Addr <=  "0001111001110";
		Trees_din <= x"4a02171c";
		wait for Clk_period;
		Addr <=  "0001111001111";
		Trees_din <= x"9400fb10";
		wait for Clk_period;
		Addr <=  "0001111010000";
		Trees_din <= x"2f022808";
		wait for Clk_period;
		Addr <=  "0001111010001";
		Trees_din <= x"c902a304";
		wait for Clk_period;
		Addr <=  "0001111010010";
		Trees_din <= x"00200fa5";
		wait for Clk_period;
		Addr <=  "0001111010011";
		Trees_din <= x"ffa70fa5";
		wait for Clk_period;
		Addr <=  "0001111010100";
		Trees_din <= x"6200d104";
		wait for Clk_period;
		Addr <=  "0001111010101";
		Trees_din <= x"ffe50fa5";
		wait for Clk_period;
		Addr <=  "0001111010110";
		Trees_din <= x"00730fa5";
		wait for Clk_period;
		Addr <=  "0001111010111";
		Trees_din <= x"65002004";
		wait for Clk_period;
		Addr <=  "0001111011000";
		Trees_din <= x"00140fa5";
		wait for Clk_period;
		Addr <=  "0001111011001";
		Trees_din <= x"ce03e904";
		wait for Clk_period;
		Addr <=  "0001111011010";
		Trees_din <= x"ff790fa5";
		wait for Clk_period;
		Addr <=  "0001111011011";
		Trees_din <= x"ffe90fa5";
		wait for Clk_period;
		Addr <=  "0001111011100";
		Trees_din <= x"8701ab10";
		wait for Clk_period;
		Addr <=  "0001111011101";
		Trees_din <= x"f500d108";
		wait for Clk_period;
		Addr <=  "0001111011110";
		Trees_din <= x"2f02f004";
		wait for Clk_period;
		Addr <=  "0001111011111";
		Trees_din <= x"ffd10fa5";
		wait for Clk_period;
		Addr <=  "0001111100000";
		Trees_din <= x"00510fa5";
		wait for Clk_period;
		Addr <=  "0001111100001";
		Trees_din <= x"a3017904";
		wait for Clk_period;
		Addr <=  "0001111100010";
		Trees_din <= x"00180fa5";
		wait for Clk_period;
		Addr <=  "0001111100011";
		Trees_din <= x"00930fa5";
		wait for Clk_period;
		Addr <=  "0001111100100";
		Trees_din <= x"be006408";
		wait for Clk_period;
		Addr <=  "0001111100101";
		Trees_din <= x"54009f04";
		wait for Clk_period;
		Addr <=  "0001111100110";
		Trees_din <= x"004e0fa5";
		wait for Clk_period;
		Addr <=  "0001111100111";
		Trees_din <= x"fff80fa5";
		wait for Clk_period;
		Addr <=  "0001111101000";
		Trees_din <= x"ffb20fa5";
		wait for Clk_period;
		Addr <=  "0001111101001";
		Trees_din <= x"2601d824";
		wait for Clk_period;
		Addr <=  "0001111101010";
		Trees_din <= x"62018710";
		wait for Clk_period;
		Addr <=  "0001111101011";
		Trees_din <= x"b802f208";
		wait for Clk_period;
		Addr <=  "0001111101100";
		Trees_din <= x"51009a04";
		wait for Clk_period;
		Addr <=  "0001111101101";
		Trees_din <= x"ffdf1009";
		wait for Clk_period;
		Addr <=  "0001111101110";
		Trees_din <= x"ff821009";
		wait for Clk_period;
		Addr <=  "0001111101111";
		Trees_din <= x"bb010d04";
		wait for Clk_period;
		Addr <=  "0001111110000";
		Trees_din <= x"00261009";
		wait for Clk_period;
		Addr <=  "0001111110001";
		Trees_din <= x"ffbe1009";
		wait for Clk_period;
		Addr <=  "0001111110010";
		Trees_din <= x"ca003908";
		wait for Clk_period;
		Addr <=  "0001111110011";
		Trees_din <= x"0c020b04";
		wait for Clk_period;
		Addr <=  "0001111110100";
		Trees_din <= x"000e1009";
		wait for Clk_period;
		Addr <=  "0001111110101";
		Trees_din <= x"00711009";
		wait for Clk_period;
		Addr <=  "0001111110110";
		Trees_din <= x"e600f108";
		wait for Clk_period;
		Addr <=  "0001111110111";
		Trees_din <= x"1402a604";
		wait for Clk_period;
		Addr <=  "0001111111000";
		Trees_din <= x"ffe81009";
		wait for Clk_period;
		Addr <=  "0001111111001";
		Trees_din <= x"00481009";
		wait for Clk_period;
		Addr <=  "0001111111010";
		Trees_din <= x"ffa91009";
		wait for Clk_period;
		Addr <=  "0001111111011";
		Trees_din <= x"41017608";
		wait for Clk_period;
		Addr <=  "0001111111100";
		Trees_din <= x"fa025704";
		wait for Clk_period;
		Addr <=  "0001111111101";
		Trees_din <= x"ffb61009";
		wait for Clk_period;
		Addr <=  "0001111111110";
		Trees_din <= x"00491009";
		wait for Clk_period;
		Addr <=  "0001111111111";
		Trees_din <= x"25020504";
		wait for Clk_period;
		Addr <=  "0010000000000";
		Trees_din <= x"00901009";
		wait for Clk_period;
		Addr <=  "0010000000001";
		Trees_din <= x"00051009";
		wait for Clk_period;
		Addr <=  "0010000000010";
		Trees_din <= x"4a02bc20";
		wait for Clk_period;
		Addr <=  "0010000000011";
		Trees_din <= x"94017a18";
		wait for Clk_period;
		Addr <=  "0010000000100";
		Trees_din <= x"30019008";
		wait for Clk_period;
		Addr <=  "0010000000101";
		Trees_din <= x"22018c04";
		wait for Clk_period;
		Addr <=  "0010000000110";
		Trees_din <= x"ffa91065";
		wait for Clk_period;
		Addr <=  "0010000000111";
		Trees_din <= x"000e1065";
		wait for Clk_period;
		Addr <=  "0010000001000";
		Trees_din <= x"c903e508";
		wait for Clk_period;
		Addr <=  "0010000001001";
		Trees_din <= x"4a011f04";
		wait for Clk_period;
		Addr <=  "0010000001010";
		Trees_din <= x"00191065";
		wait for Clk_period;
		Addr <=  "0010000001011";
		Trees_din <= x"00751065";
		wait for Clk_period;
		Addr <=  "0010000001100";
		Trees_din <= x"2f030704";
		wait for Clk_period;
		Addr <=  "0010000001101";
		Trees_din <= x"ffcd1065";
		wait for Clk_period;
		Addr <=  "0010000001110";
		Trees_din <= x"00311065";
		wait for Clk_period;
		Addr <=  "0010000001111";
		Trees_din <= x"7002a804";
		wait for Clk_period;
		Addr <=  "0010000010000";
		Trees_din <= x"ff831065";
		wait for Clk_period;
		Addr <=  "0010000010001";
		Trees_din <= x"fff11065";
		wait for Clk_period;
		Addr <=  "0010000010010";
		Trees_din <= x"eb00e608";
		wait for Clk_period;
		Addr <=  "0010000010011";
		Trees_din <= x"b601c304";
		wait for Clk_period;
		Addr <=  "0010000010100";
		Trees_din <= x"002a1065";
		wait for Clk_period;
		Addr <=  "0010000010101";
		Trees_din <= x"00911065";
		wait for Clk_period;
		Addr <=  "0010000010110";
		Trees_din <= x"99002c04";
		wait for Clk_period;
		Addr <=  "0010000010111";
		Trees_din <= x"003f1065";
		wait for Clk_period;
		Addr <=  "0010000011000";
		Trees_din <= x"ffd41065";
		wait for Clk_period;
		Addr <=  "0010000011001";
		Trees_din <= x"2601aa1c";
		wait for Clk_period;
		Addr <=  "0010000011010";
		Trees_din <= x"99000b08";
		wait for Clk_period;
		Addr <=  "0010000011011";
		Trees_din <= x"22029604";
		wait for Clk_period;
		Addr <=  "0010000011100";
		Trees_din <= x"fffa10c1";
		wait for Clk_period;
		Addr <=  "0010000011101";
		Trees_din <= x"005c10c1";
		wait for Clk_period;
		Addr <=  "0010000011110";
		Trees_din <= x"54009008";
		wait for Clk_period;
		Addr <=  "0010000011111";
		Trees_din <= x"0903a004";
		wait for Clk_period;
		Addr <=  "0010000100000";
		Trees_din <= x"ffca10c1";
		wait for Clk_period;
		Addr <=  "0010000100001";
		Trees_din <= x"003a10c1";
		wait for Clk_period;
		Addr <=  "0010000100010";
		Trees_din <= x"cb041a08";
		wait for Clk_period;
		Addr <=  "0010000100011";
		Trees_din <= x"9400d204";
		wait for Clk_period;
		Addr <=  "0010000100100";
		Trees_din <= x"ffd510c1";
		wait for Clk_period;
		Addr <=  "0010000100101";
		Trees_din <= x"ff8010c1";
		wait for Clk_period;
		Addr <=  "0010000100110";
		Trees_din <= x"fff210c1";
		wait for Clk_period;
		Addr <=  "0010000100111";
		Trees_din <= x"da023c10";
		wait for Clk_period;
		Addr <=  "0010000101000";
		Trees_din <= x"87012308";
		wait for Clk_period;
		Addr <=  "0010000101001";
		Trees_din <= x"8a01fc04";
		wait for Clk_period;
		Addr <=  "0010000101010";
		Trees_din <= x"002910c1";
		wait for Clk_period;
		Addr <=  "0010000101011";
		Trees_din <= x"009010c1";
		wait for Clk_period;
		Addr <=  "0010000101100";
		Trees_din <= x"b603b804";
		wait for Clk_period;
		Addr <=  "0010000101101";
		Trees_din <= x"ffdc10c1";
		wait for Clk_period;
		Addr <=  "0010000101110";
		Trees_din <= x"004410c1";
		wait for Clk_period;
		Addr <=  "0010000101111";
		Trees_din <= x"ffd110c1";
		wait for Clk_period;
		Addr <=  "0010000110000";
		Trees_din <= x"4a02bc1c";
		wait for Clk_period;
		Addr <=  "0010000110001";
		Trees_din <= x"6201740c";
		wait for Clk_period;
		Addr <=  "0010000110010";
		Trees_din <= x"a0001704";
		wait for Clk_period;
		Addr <=  "0010000110011";
		Trees_din <= x"0011110d";
		wait for Clk_period;
		Addr <=  "0010000110100";
		Trees_din <= x"54008c04";
		wait for Clk_period;
		Addr <=  "0010000110101";
		Trees_din <= x"ffe8110d";
		wait for Clk_period;
		Addr <=  "0010000110110";
		Trees_din <= x"ff90110d";
		wait for Clk_period;
		Addr <=  "0010000110111";
		Trees_din <= x"41017608";
		wait for Clk_period;
		Addr <=  "0010000111000";
		Trees_din <= x"29022e04";
		wait for Clk_period;
		Addr <=  "0010000111001";
		Trees_din <= x"ffb5110d";
		wait for Clk_period;
		Addr <=  "0010000111010";
		Trees_din <= x"0013110d";
		wait for Clk_period;
		Addr <=  "0010000111011";
		Trees_din <= x"53063204";
		wait for Clk_period;
		Addr <=  "0010000111100";
		Trees_din <= x"0066110d";
		wait for Clk_period;
		Addr <=  "0010000111101";
		Trees_din <= x"ffec110d";
		wait for Clk_period;
		Addr <=  "0010000111110";
		Trees_din <= x"51013f08";
		wait for Clk_period;
		Addr <=  "0010000111111";
		Trees_din <= x"77014804";
		wait for Clk_period;
		Addr <=  "0010001000000";
		Trees_din <= x"0021110d";
		wait for Clk_period;
		Addr <=  "0010001000001";
		Trees_din <= x"008b110d";
		wait for Clk_period;
		Addr <=  "0010001000010";
		Trees_din <= x"fff5110d";
		wait for Clk_period;
		Addr <=  "0010001000011";
		Trees_din <= x"3d01831c";
		wait for Clk_period;
		Addr <=  "0010001000100";
		Trees_din <= x"9400fb14";
		wait for Clk_period;
		Addr <=  "0010001000101";
		Trees_din <= x"04055f0c";
		wait for Clk_period;
		Addr <=  "0010001000110";
		Trees_din <= x"19028904";
		wait for Clk_period;
		Addr <=  "0010001000111";
		Trees_din <= x"ffee1161";
		wait for Clk_period;
		Addr <=  "0010001001000";
		Trees_din <= x"87014204";
		wait for Clk_period;
		Addr <=  "0010001001001";
		Trees_din <= x"00631161";
		wait for Clk_period;
		Addr <=  "0010001001010";
		Trees_din <= x"001a1161";
		wait for Clk_period;
		Addr <=  "0010001001011";
		Trees_din <= x"1f03aa04";
		wait for Clk_period;
		Addr <=  "0010001001100";
		Trees_din <= x"00021161";
		wait for Clk_period;
		Addr <=  "0010001001101";
		Trees_din <= x"ffb81161";
		wait for Clk_period;
		Addr <=  "0010001001110";
		Trees_din <= x"a601c804";
		wait for Clk_period;
		Addr <=  "0010001001111";
		Trees_din <= x"fff21161";
		wait for Clk_period;
		Addr <=  "0010001010000";
		Trees_din <= x"ff921161";
		wait for Clk_period;
		Addr <=  "0010001010001";
		Trees_din <= x"c800f708";
		wait for Clk_period;
		Addr <=  "0010001010010";
		Trees_din <= x"f500d104";
		wait for Clk_period;
		Addr <=  "0010001010011";
		Trees_din <= x"00011161";
		wait for Clk_period;
		Addr <=  "0010001010100";
		Trees_din <= x"00891161";
		wait for Clk_period;
		Addr <=  "0010001010101";
		Trees_din <= x"70025b04";
		wait for Clk_period;
		Addr <=  "0010001010110";
		Trees_din <= x"ffbf1161";
		wait for Clk_period;
		Addr <=  "0010001010111";
		Trees_din <= x"001e1161";
		wait for Clk_period;
		Addr <=  "0010001011000";
		Trees_din <= x"2601df1c";
		wait for Clk_period;
		Addr <=  "0010001011001";
		Trees_din <= x"6500b814";
		wait for Clk_period;
		Addr <=  "0010001011010";
		Trees_din <= x"03004e08";
		wait for Clk_period;
		Addr <=  "0010001011011";
		Trees_din <= x"e9019704";
		wait for Clk_period;
		Addr <=  "0010001011100";
		Trees_din <= x"fff711b5";
		wait for Clk_period;
		Addr <=  "0010001011101";
		Trees_din <= x"ffb311b5";
		wait for Clk_period;
		Addr <=  "0010001011110";
		Trees_din <= x"22018c08";
		wait for Clk_period;
		Addr <=  "0010001011111";
		Trees_din <= x"94009c04";
		wait for Clk_period;
		Addr <=  "0010001100000";
		Trees_din <= x"001c11b5";
		wait for Clk_period;
		Addr <=  "0010001100001";
		Trees_din <= x"ffd211b5";
		wait for Clk_period;
		Addr <=  "0010001100010";
		Trees_din <= x"005311b5";
		wait for Clk_period;
		Addr <=  "0010001100011";
		Trees_din <= x"bb008004";
		wait for Clk_period;
		Addr <=  "0010001100100";
		Trees_din <= x"ffe311b5";
		wait for Clk_period;
		Addr <=  "0010001100101";
		Trees_din <= x"ff9811b5";
		wait for Clk_period;
		Addr <=  "0010001100110";
		Trees_din <= x"41019a08";
		wait for Clk_period;
		Addr <=  "0010001100111";
		Trees_din <= x"fa025704";
		wait for Clk_period;
		Addr <=  "0010001101000";
		Trees_din <= x"ffc911b5";
		wait for Clk_period;
		Addr <=  "0010001101001";
		Trees_din <= x"003411b5";
		wait for Clk_period;
		Addr <=  "0010001101010";
		Trees_din <= x"87019e04";
		wait for Clk_period;
		Addr <=  "0010001101011";
		Trees_din <= x"008511b5";
		wait for Clk_period;
		Addr <=  "0010001101100";
		Trees_din <= x"001711b5";
		wait for Clk_period;
		Addr <=  "0010001101101";
		Trees_din <= x"0c028214";
		wait for Clk_period;
		Addr <=  "0010001101110";
		Trees_din <= x"5901620c";
		wait for Clk_period;
		Addr <=  "0010001101111";
		Trees_din <= x"64046708";
		wait for Clk_period;
		Addr <=  "0010001110000";
		Trees_din <= x"9a04a304";
		wait for Clk_period;
		Addr <=  "0010001110001";
		Trees_din <= x"ff9b11f1";
		wait for Clk_period;
		Addr <=  "0010001110010";
		Trees_din <= x"ffe611f1";
		wait for Clk_period;
		Addr <=  "0010001110011";
		Trees_din <= x"000d11f1";
		wait for Clk_period;
		Addr <=  "0010001110100";
		Trees_din <= x"93008104";
		wait for Clk_period;
		Addr <=  "0010001110101";
		Trees_din <= x"004811f1";
		wait for Clk_period;
		Addr <=  "0010001110110";
		Trees_din <= x"ffdf11f1";
		wait for Clk_period;
		Addr <=  "0010001110111";
		Trees_din <= x"a000bc08";
		wait for Clk_period;
		Addr <=  "0010001111000";
		Trees_din <= x"3d00c004";
		wait for Clk_period;
		Addr <=  "0010001111001";
		Trees_din <= x"001311f1";
		wait for Clk_period;
		Addr <=  "0010001111010";
		Trees_din <= x"007f11f1";
		wait for Clk_period;
		Addr <=  "0010001111011";
		Trees_din <= x"ffcf11f1";
		wait for Clk_period;
		Addr <=  "0010001111100";
		Trees_din <= x"f4012b14";
		wait for Clk_period;
		Addr <=  "0010001111101";
		Trees_din <= x"0c016908";
		wait for Clk_period;
		Addr <=  "0010001111110";
		Trees_din <= x"3001e604";
		wait for Clk_period;
		Addr <=  "0010001111111";
		Trees_din <= x"ffc7122d";
		wait for Clk_period;
		Addr <=  "0010010000000";
		Trees_din <= x"0017122d";
		wait for Clk_period;
		Addr <=  "0010010000001";
		Trees_din <= x"7a019508";
		wait for Clk_period;
		Addr <=  "0010010000010";
		Trees_din <= x"17021d04";
		wait for Clk_period;
		Addr <=  "0010010000011";
		Trees_din <= x"ffe6122d";
		wait for Clk_period;
		Addr <=  "0010010000100";
		Trees_din <= x"0039122d";
		wait for Clk_period;
		Addr <=  "0010010000101";
		Trees_din <= x"007c122d";
		wait for Clk_period;
		Addr <=  "0010010000110";
		Trees_din <= x"8700eb08";
		wait for Clk_period;
		Addr <=  "0010010000111";
		Trees_din <= x"e600f104";
		wait for Clk_period;
		Addr <=  "0010010001000";
		Trees_din <= x"002e122d";
		wait for Clk_period;
		Addr <=  "0010010001001";
		Trees_din <= x"ffce122d";
		wait for Clk_period;
		Addr <=  "0010010001010";
		Trees_din <= x"ff9c122d";
		wait for Clk_period;
		Addr <=  "0010010001011";
		Trees_din <= x"2501f218";
		wait for Clk_period;
		Addr <=  "0010010001100";
		Trees_din <= x"c4029b10";
		wait for Clk_period;
		Addr <=  "0010010001101";
		Trees_din <= x"1402d308";
		wait for Clk_period;
		Addr <=  "0010010001110";
		Trees_din <= x"3d018304";
		wait for Clk_period;
		Addr <=  "0010010001111";
		Trees_din <= x"ffbb1269";
		wait for Clk_period;
		Addr <=  "0010010010000";
		Trees_din <= x"00131269";
		wait for Clk_period;
		Addr <=  "0010010010001";
		Trees_din <= x"d5004a04";
		wait for Clk_period;
		Addr <=  "0010010010010";
		Trees_din <= x"00491269";
		wait for Clk_period;
		Addr <=  "0010010010011";
		Trees_din <= x"000f1269";
		wait for Clk_period;
		Addr <=  "0010010010100";
		Trees_din <= x"41017604";
		wait for Clk_period;
		Addr <=  "0010010010101";
		Trees_din <= x"000a1269";
		wait for Clk_period;
		Addr <=  "0010010010110";
		Trees_din <= x"00771269";
		wait for Clk_period;
		Addr <=  "0010010010111";
		Trees_din <= x"81009704";
		wait for Clk_period;
		Addr <=  "0010010011000";
		Trees_din <= x"00001269";
		wait for Clk_period;
		Addr <=  "0010010011001";
		Trees_din <= x"ffa81269";
		wait for Clk_period;
		Addr <=  "0010010011010";
		Trees_din <= x"5400d010";
		wait for Clk_period;
		Addr <=  "0010010011011";
		Trees_din <= x"41017608";
		wait for Clk_period;
		Addr <=  "0010010011100";
		Trees_din <= x"29022e04";
		wait for Clk_period;
		Addr <=  "0010010011101";
		Trees_din <= x"ffc8129d";
		wait for Clk_period;
		Addr <=  "0010010011110";
		Trees_din <= x"0018129d";
		wait for Clk_period;
		Addr <=  "0010010011111";
		Trees_din <= x"3700cb04";
		wait for Clk_period;
		Addr <=  "0010010100000";
		Trees_din <= x"0009129d";
		wait for Clk_period;
		Addr <=  "0010010100001";
		Trees_din <= x"0073129d";
		wait for Clk_period;
		Addr <=  "0010010100010";
		Trees_din <= x"2f02f008";
		wait for Clk_period;
		Addr <=  "0010010100011";
		Trees_din <= x"99003304";
		wait for Clk_period;
		Addr <=  "0010010100100";
		Trees_din <= x"ffed129d";
		wait for Clk_period;
		Addr <=  "0010010100101";
		Trees_din <= x"ffa3129d";
		wait for Clk_period;
		Addr <=  "0010010100110";
		Trees_din <= x"0013129d";
		wait for Clk_period;
		Addr <=  "0010010100111";
		Trees_din <= x"2f020e0c";
		wait for Clk_period;
		Addr <=  "0010010101000";
		Trees_din <= x"e0004004";
		wait for Clk_period;
		Addr <=  "0010010101001";
		Trees_din <= x"001112d1";
		wait for Clk_period;
		Addr <=  "0010010101010";
		Trees_din <= x"e600e704";
		wait for Clk_period;
		Addr <=  "0010010101011";
		Trees_din <= x"ffe712d1";
		wait for Clk_period;
		Addr <=  "0010010101100";
		Trees_din <= x"ffa412d1";
		wait for Clk_period;
		Addr <=  "0010010101101";
		Trees_din <= x"94017a0c";
		wait for Clk_period;
		Addr <=  "0010010101110";
		Trees_din <= x"0406b308";
		wait for Clk_period;
		Addr <=  "0010010101111";
		Trees_din <= x"fe014404";
		wait for Clk_period;
		Addr <=  "0010010110000";
		Trees_din <= x"001812d1";
		wait for Clk_period;
		Addr <=  "0010010110001";
		Trees_din <= x"007412d1";
		wait for Clk_period;
		Addr <=  "0010010110010";
		Trees_din <= x"fff112d1";
		wait for Clk_period;
		Addr <=  "0010010110011";
		Trees_din <= x"ffd712d1";
		wait for Clk_period;
		Addr <=  "0010010110100";
		Trees_din <= x"6201870c";
		wait for Clk_period;
		Addr <=  "0010010110101";
		Trees_din <= x"8100a108";
		wait for Clk_period;
		Addr <=  "0010010110110";
		Trees_din <= x"63002e04";
		wait for Clk_period;
		Addr <=  "0010010110111";
		Trees_din <= x"ffe01305";
		wait for Clk_period;
		Addr <=  "0010010111000";
		Trees_din <= x"00241305";
		wait for Clk_period;
		Addr <=  "0010010111001";
		Trees_din <= x"ffb31305";
		wait for Clk_period;
		Addr <=  "0010010111010";
		Trees_din <= x"4101a508";
		wait for Clk_period;
		Addr <=  "0010010111011";
		Trees_din <= x"5b026e04";
		wait for Clk_period;
		Addr <=  "0010010111100";
		Trees_din <= x"ffd11305";
		wait for Clk_period;
		Addr <=  "0010010111101";
		Trees_din <= x"00141305";
		wait for Clk_period;
		Addr <=  "0010010111110";
		Trees_din <= x"5c01ae04";
		wait for Clk_period;
		Addr <=  "0010010111111";
		Trees_din <= x"00071305";
		wait for Clk_period;
		Addr <=  "0010011000000";
		Trees_din <= x"006c1305";
		wait for Clk_period;
		Addr <=  "0010011000001";
		Trees_din <= x"c001f314";
		wait for Clk_period;
		Addr <=  "0010011000010";
		Trees_din <= x"2f02f00c";
		wait for Clk_period;
		Addr <=  "0010011000011";
		Trees_din <= x"4101b804";
		wait for Clk_period;
		Addr <=  "0010011000100";
		Trees_din <= x"ffca1339";
		wait for Clk_period;
		Addr <=  "0010011000101";
		Trees_din <= x"5400b104";
		wait for Clk_period;
		Addr <=  "0010011000110";
		Trees_din <= x"003c1339";
		wait for Clk_period;
		Addr <=  "0010011000111";
		Trees_din <= x"ffed1339";
		wait for Clk_period;
		Addr <=  "0010011001000";
		Trees_din <= x"16007204";
		wait for Clk_period;
		Addr <=  "0010011001001";
		Trees_din <= x"00071339";
		wait for Clk_period;
		Addr <=  "0010011001010";
		Trees_din <= x"006e1339";
		wait for Clk_period;
		Addr <=  "0010011001011";
		Trees_din <= x"19048604";
		wait for Clk_period;
		Addr <=  "0010011001100";
		Trees_din <= x"ffae1339";
		wait for Clk_period;
		Addr <=  "0010011001101";
		Trees_din <= x"fff61339";
		wait for Clk_period;
		Addr <=  "0010011001110";
		Trees_din <= x"f4012b10";
		wait for Clk_period;
		Addr <=  "0010011001111";
		Trees_din <= x"29023e08";
		wait for Clk_period;
		Addr <=  "0010011010000";
		Trees_din <= x"c7010b04";
		wait for Clk_period;
		Addr <=  "0010011010001";
		Trees_din <= x"ffd01365";
		wait for Clk_period;
		Addr <=  "0010011010010";
		Trees_din <= x"00161365";
		wait for Clk_period;
		Addr <=  "0010011010011";
		Trees_din <= x"87010504";
		wait for Clk_period;
		Addr <=  "0010011010100";
		Trees_din <= x"006a1365";
		wait for Clk_period;
		Addr <=  "0010011010101";
		Trees_din <= x"000a1365";
		wait for Clk_period;
		Addr <=  "0010011010110";
		Trees_din <= x"8700eb04";
		wait for Clk_period;
		Addr <=  "0010011010111";
		Trees_din <= x"fffb1365";
		wait for Clk_period;
		Addr <=  "0010011011000";
		Trees_din <= x"ffae1365";
		wait for Clk_period;
		Addr <=  "0010011011001";
		Trees_din <= x"eb008508";
		wait for Clk_period;
		Addr <=  "0010011011010";
		Trees_din <= x"5b017d04";
		wait for Clk_period;
		Addr <=  "0010011011011";
		Trees_din <= x"fff31389";
		wait for Clk_period;
		Addr <=  "0010011011100";
		Trees_din <= x"005d1389";
		wait for Clk_period;
		Addr <=  "0010011011101";
		Trees_din <= x"6101e908";
		wait for Clk_period;
		Addr <=  "0010011011110";
		Trees_din <= x"5a015604";
		wait for Clk_period;
		Addr <=  "0010011011111";
		Trees_din <= x"ffdc1389";
		wait for Clk_period;
		Addr <=  "0010011100000";
		Trees_din <= x"00271389";
		wait for Clk_period;
		Addr <=  "0010011100001";
		Trees_din <= x"ffb91389";
		wait for Clk_period;
		Addr <=  "0010011100010";
		Trees_din <= x"3d018310";
		wait for Clk_period;
		Addr <=  "0010011100011";
		Trees_din <= x"9a048f08";
		wait for Clk_period;
		Addr <=  "0010011100100";
		Trees_din <= x"a0003604";
		wait for Clk_period;
		Addr <=  "0010011100101";
		Trees_din <= x"fff613b5";
		wait for Clk_period;
		Addr <=  "0010011100110";
		Trees_din <= x"ffb313b5";
		wait for Clk_period;
		Addr <=  "0010011100111";
		Trees_din <= x"b201a904";
		wait for Clk_period;
		Addr <=  "0010011101000";
		Trees_din <= x"fff013b5";
		wait for Clk_period;
		Addr <=  "0010011101001";
		Trees_din <= x"002413b5";
		wait for Clk_period;
		Addr <=  "0010011101010";
		Trees_din <= x"b3016604";
		wait for Clk_period;
		Addr <=  "0010011101011";
		Trees_din <= x"ffe513b5";
		wait for Clk_period;
		Addr <=  "0010011101100";
		Trees_din <= x"005513b5";
		wait for Clk_period;
		Addr <=  "0010011101101";
		Trees_din <= x"62012808";
		wait for Clk_period;
		Addr <=  "0010011101110";
		Trees_din <= x"81009204";
		wait for Clk_period;
		Addr <=  "0010011101111";
		Trees_din <= x"000113e1";
		wait for Clk_period;
		Addr <=  "0010011110000";
		Trees_din <= x"ffb713e1";
		wait for Clk_period;
		Addr <=  "0010011110001";
		Trees_din <= x"f4012b0c";
		wait for Clk_period;
		Addr <=  "0010011110010";
		Trees_din <= x"30020804";
		wait for Clk_period;
		Addr <=  "0010011110011";
		Trees_din <= x"fffd13e1";
		wait for Clk_period;
		Addr <=  "0010011110100";
		Trees_din <= x"77019304";
		wait for Clk_period;
		Addr <=  "0010011110101";
		Trees_din <= x"001513e1";
		wait for Clk_period;
		Addr <=  "0010011110110";
		Trees_din <= x"005e13e1";
		wait for Clk_period;
		Addr <=  "0010011110111";
		Trees_din <= x"ffe713e1";
		wait for Clk_period;
		Addr <=  "0010011111000";
		Trees_din <= x"2f02f00c";
		wait for Clk_period;
		Addr <=  "0010011111001";
		Trees_din <= x"99000f04";
		wait for Clk_period;
		Addr <=  "0010011111010";
		Trees_din <= x"00181405";
		wait for Clk_period;
		Addr <=  "0010011111011";
		Trees_din <= x"59017004";
		wait for Clk_period;
		Addr <=  "0010011111100";
		Trees_din <= x"ffb71405";
		wait for Clk_period;
		Addr <=  "0010011111101";
		Trees_din <= x"fffc1405";
		wait for Clk_period;
		Addr <=  "0010011111110";
		Trees_din <= x"bb012b04";
		wait for Clk_period;
		Addr <=  "0010011111111";
		Trees_din <= x"004f1405";
		wait for Clk_period;
		Addr <=  "0010100000000";
		Trees_din <= x"fff11405";
		wait for Clk_period;
		Addr <=  "0010100000001";
		Trees_din <= x"ca008910";
		wait for Clk_period;
		Addr <=  "0010100000010";
		Trees_din <= x"5c01c508";
		wait for Clk_period;
		Addr <=  "0010100000011";
		Trees_din <= x"f4008704";
		wait for Clk_period;
		Addr <=  "0010100000100";
		Trees_din <= x"00141431";
		wait for Clk_period;
		Addr <=  "0010100000101";
		Trees_din <= x"ffd71431";
		wait for Clk_period;
		Addr <=  "0010100000110";
		Trees_din <= x"3d016504";
		wait for Clk_period;
		Addr <=  "0010100000111";
		Trees_din <= x"00111431";
		wait for Clk_period;
		Addr <=  "0010100001000";
		Trees_din <= x"00571431";
		wait for Clk_period;
		Addr <=  "0010100001001";
		Trees_din <= x"25014704";
		wait for Clk_period;
		Addr <=  "0010100001010";
		Trees_din <= x"fffe1431";
		wait for Clk_period;
		Addr <=  "0010100001011";
		Trees_din <= x"ffbc1431";
		wait for Clk_period;
		Addr <=  "0010100001100";
		Trees_din <= x"65011410";
		wait for Clk_period;
		Addr <=  "0010100001101";
		Trees_din <= x"0c02d90c";
		wait for Clk_period;
		Addr <=  "0010100001110";
		Trees_din <= x"14031a08";
		wait for Clk_period;
		Addr <=  "0010100001111";
		Trees_din <= x"9601d304";
		wait for Clk_period;
		Addr <=  "0010100010000";
		Trees_din <= x"ffc71455";
		wait for Clk_period;
		Addr <=  "0010100010001";
		Trees_din <= x"00011455";
		wait for Clk_period;
		Addr <=  "0010100010010";
		Trees_din <= x"00251455";
		wait for Clk_period;
		Addr <=  "0010100010011";
		Trees_din <= x"004b1455";
		wait for Clk_period;
		Addr <=  "0010100010100";
		Trees_din <= x"ffc21455";
		wait for Clk_period;
		Addr <=  "0010100010101";
		Trees_din <= x"5400d00c";
		wait for Clk_period;
		Addr <=  "0010100010110";
		Trees_din <= x"41017604";
		wait for Clk_period;
		Addr <=  "0010100010111";
		Trees_din <= x"ffed1479";
		wait for Clk_period;
		Addr <=  "0010100011000";
		Trees_din <= x"92038c04";
		wait for Clk_period;
		Addr <=  "0010100011001";
		Trees_din <= x"00161479";
		wait for Clk_period;
		Addr <=  "0010100011010";
		Trees_din <= x"00531479";
		wait for Clk_period;
		Addr <=  "0010100011011";
		Trees_din <= x"99003b04";
		wait for Clk_period;
		Addr <=  "0010100011100";
		Trees_din <= x"00071479";
		wait for Clk_period;
		Addr <=  "0010100011101";
		Trees_din <= x"ffc31479";
		wait for Clk_period;
		Addr <=  "0010100011110";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  2
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"320a593c";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"0009512c";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"400c531c";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"0006b00c";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"bc0e6208";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"8c0ab704";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"ff4e00cd";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"ffbb00cd";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"001200cd";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"5e018e08";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"6a021404";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"028000cd";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"ff7800cd";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"2d0c4404";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"ff5500cd";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"002700cd";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"1b00e008";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"0e047a04";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"02a700cd";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"00b200cd";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"1100ef04";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"002700cd";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"ff5f00cd";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"78026d08";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"4d059e04";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"03b200cd";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"fff100cd";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"83080104";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"ff5b00cd";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"013c00cd";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"8c04aa18";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"5d02570c";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"5a070004";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"030800cd";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"0201e604";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"ff8100cd";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"002700cd";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"cc08cf08";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"41097104";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"ff5300cd";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"002700cd";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"01c600cd";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"78063110";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"c603c508";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"00047d04";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"ff8f00cd";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"018700cd";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"57086504";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"041f00cd";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"015400cd";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"ff6400cd";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"32091c38";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"00095124";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"400c5318";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"8c07bc0c";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"bc0e6208";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"0007eb04";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"ff550179";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"ffb20179";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"00170179";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"df00ad08";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"10067404";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"ff9c0179";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"01cc0179";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"ff620179";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"1b00e008";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"45036104";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"01c00179";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"00290179";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"ff640179";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"5e043f0c";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"37011604";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"ff8f0179";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"f6061a04";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"01c10179";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"00910179";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"5f063604";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"ff650179";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"00350179";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"0001eb0c";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"600f8b04";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"ff570179";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"47096604";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"01760179";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"ff890179";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"1a0acd10";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"04015904";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"ff850179";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"a8127d08";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"44094e04";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"01b50179";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"001b0179";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"ff900179";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"ff680179";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"3206f334";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"400d4d28";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"2d089318";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"f6001708";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"60005904";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"003d0235";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"ff960235";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"100c4e08";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"9b0f0204";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"ff580235";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"ff980235";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"7f004f04";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"ff7c0235";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"002f0235";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"6a023808";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"0a012b04";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"01350235";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"00240235";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"18001c04";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"00420235";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"ff5f0235";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"0003e404";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"ff730235";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"0300e204";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"01200235";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"00610235";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"8c028f10";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"350ce10c";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"3214f608";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"4109b604";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"ff5b0235";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"002c0235";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"00620235";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"01180235";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"1002df08";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"4018dc04";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"ff620235";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"00850235";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"44094e0c";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"78063108";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"110b5904";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"01380235";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"ff9c0235";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"ff960235";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"00088e04";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"ff750235";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"00d40235";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"3206f330";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"400d4d28";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"2d089318";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"f6001708";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"f1011c04";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"003b02f1";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"ff9e02f1";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"100c4e08";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"9b0f0204";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"ff5c02f1";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"ffa302f1";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"5b047b04";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"ff8302f1";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"002902f1";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"6a023808";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"0a012b04";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"00fc02f1";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"001f02f1";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"18001c04";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"004302f1";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"ff6402f1";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"0003e404";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"ff7a02f1";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"00ce02f1";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"00029c14";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"4d02060c";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"6c05f704";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"ff7402f1";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"8b058504";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"00f202f1";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"fff002f1";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"84161704";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"ff5f02f1";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"002d02f1";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"1002c708";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"a504ff04";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"ff6c02f1";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"007902f1";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"4f08350c";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"04011e04";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"ff9602f1";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"78063104";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"010002f1";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"ffe502f1";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"3f004c04";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"001002f1";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"ff8802f1";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"3206f324";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"400d4d18";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"2d08930c";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"0006b004";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"ff5e038d";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"c9076604";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"ff6a038d";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"00bb038d";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"6f039108";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"0f00c504";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"0076038d";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"ff67038d";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"00c8038d";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"0003e404";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"ff81038d";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"3202ad04";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"0020038d";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"00c3038d";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"00029c14";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"600cf908";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"a6046104";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"002d038d";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"ff63038d";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"47096608";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"4d043d04";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"00d2038d";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"ffac038d";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"ff82038d";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"1a0acd14";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"04013204";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"ff8e038d";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"55091b08";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"8b0ef504";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"00dc038d";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"ffc5038d";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"160c1a04";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"ff88038d";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"004f038d";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"ff76038d";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"3206f328";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"400d4d1c";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"2d08930c";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"0006b004";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"ff600451";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"c9076604";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"ff6f0451";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"009f0451";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"5b063508";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"b5030d04";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"ff6d0451";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"fff60451";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"5701f604";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"00ff0451";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"ffa40451";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"0003e404";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"ff880451";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"1b00eb04";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"00ae0451";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"002e0451";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"0003261c";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"600d8f0c";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"2f01b704";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"ff640451";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"48066b04";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"ffaa0451";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"00830451";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"c6048a04";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"ff920451";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"2b024404";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"ffe30451";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"7101c704";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"00cc0451";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"00420451";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"1002c708";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"76029604";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"004c0451";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"ff780451";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"4f06e010";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"7e00cd08";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"44017204";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"00980451";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"ff810451";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"2200a204";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"002e0451";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"00cd0451";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"d401c804";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"00390451";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"ff920451";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"3206f324";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"400d4d18";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"2d04f704";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"ff6204f5";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"b2036708";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"8f013304";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"003904f5";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"ff6704f5";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"1902e904";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"ffa304f5";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"70010104";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"00ef04f5";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"003004f5";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"0003e404";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"ff9004f5";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"d703d004";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"002404f5";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"009a04f5";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"8c028f10";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"35032204";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"ff6b04f5";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"5304c004";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"ff9204f5";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"2d09a204";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"ffeb04f5";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"00b704f5";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"1002df08";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"8604c604";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"ff7b04f5";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"003704f5";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"2200c408";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"320f5a04";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"ff7d04f5";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"006b04f5";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"b007a008";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"27049004";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"ffe004f5";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"00bb04f5";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"b201b504";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"ff9e04f5";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"007a04f5";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"3206f328";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"00067218";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"670bee10";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"ab001608";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"ad004804";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"0065059d";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"ff87059d";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"8c0ab704";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"ff63059d";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"fffb059d";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"dd0a9004";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"ffa1059d";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"008a059d";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"41006108";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"b2013b04";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"ffab059d";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"00ab059d";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"53061f04";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"ff78059d";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"ffe8059d";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"00032614";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"600d8f08";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"2f01b704";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"ff6c059d";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"0020059d";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"cc022808";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"b5000604";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"0037059d";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"ff99059d";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"0098059d";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"55091b10";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"04015304";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"ffa3059d";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"4d0a8608";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"78060a04";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"00af059d";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"ffe5059d";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"ffca059d";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"37051b04";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"ff88059d";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"0005059d";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"3206901c";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"00067210";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"96000008";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"b202f604";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"ff970631";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"00660631";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"f1110404";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"ff640631";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"ffed0631";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"41013508";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"5d01b604";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"00950631";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"ffa90631";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"ff7e0631";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"00025e10";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"600f8b08";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"8c05f404";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"ff710631";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"000a0631";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"7101c704";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"00720631";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"ffcf0631";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"1a09681c";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"44078910";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"a8105f08";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"2704c804";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"fff10631";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"00a90631";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"2b09f504";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"ffa60631";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"00310631";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"600cf908";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"a6084c04";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"00170631";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"ff7a0631";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"00850631";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"ff9b0631";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"27056510";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"00055404";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"ff6506ad";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"ed064f04";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"ff7c06ad";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"7101dd04";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"007106ad";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"001a06ad";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"1005f214";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"5d03420c";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"55046608";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"aa021e04";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"000606ad";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"009006ad";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"ffa606ad";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"7e081204";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"ff7006ad";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"001806ad";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"44078910";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"c3002f04";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"ffff06ad";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"2d046504";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"ffff06ad";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"18060804";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"00a606ad";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"001906ad";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"00064104";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"ff8306ad";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"100c4e04";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"ffc506ad";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"007e06ad";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"3206901c";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"00067210";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"96000008";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"7e02c004";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"ffac0741";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"00410741";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"f1110404";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"ff660741";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"fff80741";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"2905d804";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"ff950741";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"6401d804";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"007b0741";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"ffee0741";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"00059e1c";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"44062a14";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"6008ad08";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"a7035c04";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"ff920741";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"001b0741";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"8907c308";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"04027904";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"00180741";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"00940741";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"ffdb0741";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"4600c504";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"00140741";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"ff750741";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"1a096810";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"45091a08";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"60059b04";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"00240741";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"00a10741";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"5d013e04";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"00550741";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"ffce0741";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"ffb30741";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"27056510";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"00055404";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"ff6707b5";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"ed052504";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"ff8307b5";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"fb023104";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"001007b5";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"005a07b5";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"10049110";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"dd085e08";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"7e042004";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"ff7b07b5";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"ffdf07b5";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"c7063a04";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"ffdb07b5";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"006d07b5";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"5a05d410";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"ab06230c";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"2d046504";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"000107b5";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"6b01b004";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"002307b5";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"009c07b5";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"ffef07b5";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"100e1308";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"9c017e04";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"ff8407b5";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"001607b5";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"006f07b5";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"32069018";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"0006720c";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"3c000304";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"fffc0831";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"96000004";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"ffe40831";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"ff670831";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"2905d804";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"ffa40831";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"59016804";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"00660831";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"00030831";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"00059e18";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"4404250c";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"6008ad04";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"ffc30831";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"4902e104";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"007d0831";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"ffff0831";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"6011f308";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"7b01e804";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"ff7d0831";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"ffe00831";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"00330831";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"5e07a20c";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"45091a08";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"1a053504";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"009a0831";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"00320831";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"00150831";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"ffc60831";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"2705650c";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"00055404";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"ff690895";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"ed052504";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"ff900895";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"003d0895";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"7e02e814";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"5d03a60c";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"5a065908";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"0804a904";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"00040895";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"007a0895";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"ffbf0895";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"600e0a04";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"ff7f0895";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"fffb0895";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"c6038108";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"e4021704";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"ffa70895";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"00190895";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"8c02f704";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"fffb0895";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"55057c04";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"00950895";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"00250895";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"2d075a10";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"00067208";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"ab001604";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"ffef08f1";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"ff6a08f1";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"5e02f504";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"004c08f1";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"ffac08f1";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"4d059e18";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"04028308";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"c302d204";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"ffab08f1";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"003208f1";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"4409240c";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"3107d408";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"2d083a04";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"002a08f1";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"009408f1";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"001508f1";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"ffea08f1";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"840e2904";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"ff9408f1";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"003d08f1";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"2705650c";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"00055404";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"ff6b0949";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"ed064f04";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"ffa20949";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"00370949";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"0005d514";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"1105020c";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"44062a08";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"f5008704";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"00750949";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"fff50949";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"ffc60949";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"400c5304";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"ff890949";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"fff50949";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"10049104";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"ffdb0949";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"04031404";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"00120949";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"008e0949";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"2d075a10";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"00067208";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"e20b7004";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"ff6d099d";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"ffe4099d";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"c6055c04";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"ffb1099d";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"003b099d";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"8907c310";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"48015204";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"ffed099d";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"8c019d04";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"0001099d";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"43016604";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"002c099d";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"008f099d";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"320f5a08";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"4005e404";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"ff95099d";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"0002099d";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"0048099d";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"27056508";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"00055404";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"ff6e09e9";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"ffe209e9";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"5d05da14";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"1b038710";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"00030908";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"1302ee04";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"003c09e9";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"ffe109e9";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"2d06c604";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"002409e9";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"008909e9";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"ffd309e9";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"2d0ab204";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"ff9d09e9";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"4402bb04";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"004809e9";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"ffe509e9";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"2d041604";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"ff710a25";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"00053210";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"44042508";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"1c014604";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"004b0a25";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"ffdc0a25";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"1800be04";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"fff20a25";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"ff920a25";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"a80b3a08";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"04031404";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"00150a25";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"00850a25";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"ffe30a25";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"3204fc08";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"8408a404";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"ff740a59";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"ffef0a59";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"5503ab0c";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"c604c804";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"ffe30a59";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"8c028504";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"00130a59";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"007d0a59";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"5d020004";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"00320a59";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"ffab0a59";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"2d08930c";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"4008a708";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"0006b004";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"ff770a8d";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"ffe20a8d";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"000f0a8d";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"89080b08";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"0f06bc04";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"00780a8d";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"00100a8d";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"320e5c04";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"ffb50a8d";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"00320a8d";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"bf074d0c";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"0006b008";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"2d05b604";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"ff780ac1";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"ffd60ac1";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"fffd0ac1";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"4409240c";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"1005f204";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"fff80ac1";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"b005ad04";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"007c0ac1";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"00190ac1";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"ffbc0ac1";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"10049108";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"8508fc04";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"ff7e0aed";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"fff20aed";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"0004c308";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"48058804";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"ffa90aed";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"001a0aed";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"5503c704";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"00740aed";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"000c0aed";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"bf074d08";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"3206f304";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"ff880b19";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"fffa0b19";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"11044d08";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"0003ab04";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"00120b19";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"006c0b19";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"8905c604";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"00290b19";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"ffbe0b19";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"10049108";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"dd07d204";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"ff880b45";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"ffea0b45";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"0004c308";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"ab008204";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"00240b45";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"ffbc0b45";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"b0045104";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"00680b45";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"00080b45";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"60066008";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"2d04ba04";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"ff8a0b69";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"ffe90b69";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"2202f204";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"ffd80b69";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"04038c04";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"fff50b69";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"00620b69";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"2d0ab20c";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"98064504";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"ff910b8d";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"1b015b04";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"00320b8d";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"ffcd0b8d";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"44052304";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"005c0b8d";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"fffb0b8d";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"bf074d08";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"2d04f704";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"ff960bb1";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"ffef0bb1";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"11044d08";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"44044604";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"005d0bb1";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"00150bb1";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"ffeb0bb1";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"00059e0c";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"1c004b04";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"00140bd5";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"6c05f704";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"ff960bd5";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"ffe40bd5";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"7e038604";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"fffa0bd5";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"00540bd5";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"10049104";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"ffab0bf1";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"22040704";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"ffdf0bf1";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"6c055104";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"00090bf1";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"00580bf1";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"27056504";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"ffac0c0d";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"5d026404";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"004a0c0d";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"7e02fa04";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"ffcb0c0d";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"00120c0d";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"320a5908";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"00053204";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"ffae0c29";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"00070c29";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"89055404";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"004c0c29";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"00040c29";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"600b840c";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"00067208";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"e204b504";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"ffa70c4d";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"ffeb0c4d";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"000f0c4d";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"89052604";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"00460c4d";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"000f0c4d";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"10075908";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"bc052e04";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"ffb20c69";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"00060c69";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"4f013c04";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"00450c69";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"fff80c69";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"bf074d04";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"ffc50c7d";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"5a05d404";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"00400c7d";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"ffeb0c7d";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"22040704";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"ffc90c91";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"6c055104";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"ffef0c91";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"00460c91";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"7e02e804";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"ffcc0ca5";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"4f014404";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"003f0ca5";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"fff50ca5";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"00059e08";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"1c013a04";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"00070cb9";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"ffb90cb9";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"002e0cb9";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"2d0ab208";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"98064504";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"ffba0ccd";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"00050ccd";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"002c0ccd";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"5d026404";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"00260cd9";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"ffd40cd9";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"100bb008";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"0404dc04";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"ffc40ced";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"00040ced";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"00320ced";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"4803c504";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"ffd50cf9";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"00230cf9";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  3
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"3f0fe350";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"200a272c";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"470af418";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"01144410";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"4c009208";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"0f030904";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"003100d5";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"ff5c00d5";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"140d2704";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"ff4f00d5";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"ffe000d5";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"47056a04";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"ff7a00d5";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"01c600d5";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"05034e10";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"3f063408";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"00017604";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"002700d5";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"ff8100d5";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"d2062804";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"031a00d5";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"002700d5";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"ff5d00d5";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"0402550c";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"7c026b04";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"ff8900d5";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"03036904";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"03e300d5";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"010b00d5";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"1006a910";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"5008b308";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"02013a04";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"002700d5";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"ff7500d5";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"98091904";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"032700d5";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"001200d5";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"24083504";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"ff5500d5";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"002700d5";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"20056c08";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"04014e04";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"013c00d5";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"ff6300d5";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"b904fd04";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"ff8f00d5";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"04083c0c";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"31006104";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"00e200d5";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"95008104";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"013c00d5";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"041200d5";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"007100d5";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"4708db4c";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"20080028";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"3f10ea20";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"1407b110";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"5c0b5a08";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"80000404";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"ffc201c1";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"ff5501c1";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"8eff4704";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"00ca01c1";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"ff6b01c1";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"9c00ad08";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"33021904";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"01e001c1";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"ff6e01c1";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"0a000004";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"003f01c1";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"ff5801c1";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"07057d04";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"ff7801c1";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"016201c1";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"c3006c10";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"02062d0c";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"7c027604";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"ff9501c1";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"23072504";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"01e801c1";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"fff301c1";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"ff7f01c1";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"cf00ef0c";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"68010704";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"ff7001c1";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"2f008f04";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"01a201c1";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"ff9901c1";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"910f1604";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"ff5801c1";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"009101c1";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"3f093714";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"04028d0c";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"2f015308";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"7a022604";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"000201c1";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"01e001c1";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"ff7f01c1";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"5610f504";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"ff5c01c1";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"005a01c1";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"0f0c2c10";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"100e130c";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"5b03ad08";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"8900e404";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"001a01c1";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"01c201c1";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"ff9e01c1";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"ff8d01c1";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"68030804";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"ff6e01c1";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"011f01c1";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"2008d140";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"3f0fe330";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"470af420";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"50052110";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"bd000608";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"3800cb04";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"00d40285";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"ff7a0285";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"560f4d04";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"ff590285";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"ffcf0285";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"3500a508";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"d9017004";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"016b0285";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"ff8e0285";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"af0b2604";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"ff620285";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"fff70285";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"6c02e408";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"09022304";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"011b0285";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"ffa10285";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"d607ab04";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"ff680285";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"00290285";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"0701d004";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"ff720285";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"04037608";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"25067e04";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"005c0285";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"01450285";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"fff80285";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"3f069c10";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"7c0da308";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"9c000004";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"006c0285";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"ff5d0285";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"1f052504";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"01090285";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"00240285";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"100e1310";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"0305c70c";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"7c026b04";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"ff900285";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"80060e04";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"013e0285";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"ff900285";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"ff880285";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"ff710285";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"20080044";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"3f0fe334";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"1407b11c";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"470af410";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"ae000008";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"5b003a04";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"00be0371";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"ff6e0371";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"a50b5b04";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"ff5e0371";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"ffd00371";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"63036808";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"3f063404";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"ffa40371";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"00dc0371";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"ff740371";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"2004f108";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"a9000704";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"00a30371";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"ff610371";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"6a06df08";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"470bda04";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"ff750371";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"00b80371";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"02020204";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"019d0371";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"00690371";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"0701d004";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"ff7a0371";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"9f022b08";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"23060b04";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"01070371";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"00550371";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"ffe60371";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"3f069c14";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"7c0a7408";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"dd000204";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"001a0371";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"ff610371";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"9203b408";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"bd021f04";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"ff940371";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"001c0371";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"01230371";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"c3035514";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"0305c710";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"7f01ad08";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"d402af04";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"004d0371";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"01060371";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"5e01af04";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"000f0371";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"ffa90371";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"ff840371";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"3108c208";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"a9041704";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"ff6b0371";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"00180371";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"00b50371";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"20079d3c";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"3f0fe32c";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"1407b118";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"470c9110";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"c3000008";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"6c00fd04";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"00c1044d";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"ff6d044d";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"91124204";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"ff60044d";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"fff5044d";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"2a058c04";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"ff88044d";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"009d044d";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"2004f108";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"a9000704";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"008b044d";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"ff65044d";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"fb01e508";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"2b026904";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"0114044d";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"ffa7044d";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"ff85044d";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"0701d004";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"ff82044d";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"9f022b08";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"e304f404";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"00df044d";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"0043044d";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"ffe9044d";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"7c050710";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"3c062e08";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"1e000004";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"0009044d";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"ff63044d";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"6c02f804";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"00d7044d";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"ff8e044d";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"100e1320";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"16036910";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"56044208";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"99108604";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"ff72044d";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"0009044d";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"ae026204";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"00b4044d";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"ffa0044d";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"5b028008";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"e5001c04";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"fff9044d";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"00e6044d";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"5d02e104";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"007e044d";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"ff85044d";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"ff79044d";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"20079d44";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"4708db30";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"1407b11c";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"c300000c";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"2003f304";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"ff750519";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"0701df04";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"ffaa0519";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"00f80519";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"8efab308";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"3c054704";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"ff780519";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"00df0519";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"91124204";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"ff620519";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"fffc0519";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"6a052e08";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"15001d04";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"fff90519";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"ff6b0519";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"33021908";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"2f01ef04";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"00f70519";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"ffad0519";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"ff7f0519";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"04028d0c";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"2600d908";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"a8088504";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"00da0519";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"00320519";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"ffa90519";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"220c7e04";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"ff720519";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"00410519";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"0103b00c";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"c3000904";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"00650519";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"cf008804";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"00070519";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"ff670519";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"52016610";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"0307390c";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"100e1308";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"09046a04";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"00c40519";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"ffc20519";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"ff940519";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"ff8b0519";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"3c0aaf04";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"ff700519";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"00830519";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"50081844";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"a9000e10";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"14075408";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"0602bf04";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"ff830605";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"002b0605";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"94083b04";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"00cf0605";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"000e0605";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"4c00921c";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"0703fa0c";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"850c0108";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"0400b204";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"ffe60605";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"ff660605";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"00930605";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"8203dc08";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"6e01cc04";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"ff8d0605";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"fffa0605";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"d703dd04";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"00ce0605";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"00000605";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"90000008";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"6c01c504";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"00b00605";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"ff790605";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"aa000308";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"05020a04";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"006c0605";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"ff9e0605";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"8efab304";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"ffae0605";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"ff620605";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"0406b320";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"0103760c";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"1803f304";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"ff720605";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"63026d04";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"00cb0605";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"00000605";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"20040708";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"c4031004";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"ff840605";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"00480605";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"100e1308";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"240cdb04";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"00bf0605";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"ffe10605";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"ffa90605";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"310ef310";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"140af708";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"41054e04";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"ff670605";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"ffd60605";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"010a7204";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"ffab0605";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"00890605";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"00830605";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"50081840";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"4c009220";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"0f04ab14";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"39062b08";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"4b023204";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"000406fd";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"ff8306fd";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"56014904";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"ffae06fd";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"5003be04";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"002806fd";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"00d006fd";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"a40dfb08";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"8208a904";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"ff6a06fd";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"ffde06fd";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"002a06fd";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"a9000708";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"14068d04";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"ff9a06fd";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"008c06fd";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"90000008";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"6c01c504";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"009b06fd";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"ff7f06fd";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"aa000308";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"2004b104";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"ffa606fd";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"005c06fd";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"b0003604";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"ffbe06fd";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"ff6306fd";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"0404871c";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"20040708";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"3f0d8d04";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"ff8206fd";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"003806fd";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"01036508";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"6d000804";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"006c06fd";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"ff9906fd";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"02067b08";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"bd095304";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"00b806fd";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"001306fd";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"fffd06fd";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"2b01b714";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"c9054c0c";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"08028d04";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"001706fd";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"35024a04";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"00c106fd";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"003406fd";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"8a015a04";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"ff9906fd";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"000406fd";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"0111e408";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"8d000004";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"ffd506fd";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"ff6806fd";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"003b06fd";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"50081838";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"fb00a71c";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"3e02c304";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"ff6d07c1";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"4705c00c";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"84000004";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"008707c1";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"5c081804";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"ff7807c1";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"001407c1";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"510a8708";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"cd026d04";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"fffa07c1";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"00bd07c1";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"ffef07c1";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"a9000e08";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"72005204";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"007007c1";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"ffa007c1";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"8efab308";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"f6076a04";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"ff8f07c1";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"00d507c1";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"470a4504";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"ff6507c1";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"2d01a204";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"003907c1";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"ff9807c1";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"0406b31c";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"39053f08";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"1308db04";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"ff8607c1";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"006407c1";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"02067b0c";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"0a084308";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"82014f04";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"000c07c1";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"00a907c1";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"ffc507c1";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"0f020404";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"003a07c1";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"ff9807c1";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"4c00330c";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"200b4a04";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"ffa007c1";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"c3002f04";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"008c07c1";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"fffe07c1";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"ff7407c1";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"50081838";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"4c00921c";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"0f04ab14";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"39062b08";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"59023a04";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"ff95088d";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"fff8088d";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"54027d04";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"ffee088d";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"70039004";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"00b3088d";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"002d088d";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"ce06ea04";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"ff76088d";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"0011088d";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"8efab308";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"b0012904";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"00d0088d";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"ff93088d";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"a9000708";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"1405d104";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"ffac088d";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"006a088d";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"3a000104";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"0014088d";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"b90b8f04";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"ff65088d";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"ffc1088d";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"0404871c";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"20040708";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"e504e504";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"ff92088d";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"0011088d";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"3c036408";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"0d02fa04";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"ffa8088d";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"0065088d";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"3f04a304";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"fff8088d";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"7f010504";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"00a8088d";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"002c088d";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"2b01b70c";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"3e064b04";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"ffb3088d";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"92039104";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"001a088d";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"009f088d";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"dc104504";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"ff74088d";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"000d088d";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"3905e120";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"8efab308";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"7e009d04";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"00c20939";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"ff9d0939";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"0109e40c";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"200ab604";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"ff660939";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"1306e904";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"ffa40939";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"003e0939";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"fd04a204";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"ff900939";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"81093204";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"00750939";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"ffea0939";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"16037c20";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"1f03650c";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"b9069c04";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"ff9b0939";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"0e056204";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"00aa0939";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"ffe40939";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"14072e08";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"04009c04";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"ffe50939";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"ff6d0939";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"33021908";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"3c046e04";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"001b0939";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"00640939";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"ffae0939";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"100e1314";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"2002f904";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"ffa30939";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"5b028708";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"b9022904";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"fffd0939";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"00990939";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"05012704";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"00550939";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"ffb10939";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"ff950939";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"3905e11c";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"8efab308";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"a7010d04";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"00b009dd";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"ffa409dd";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"0109e408";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"460d7904";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"ff6709dd";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"000509dd";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"fd04a204";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"ff9809dd";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"81093204";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"006a09dd";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"ffef09dd";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"16037c1c";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"1f03650c";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"b9069c04";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"ffa309dd";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"a3007804";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"ffe209dd";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"009609dd";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"14072e08";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"ce055f04";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"ff7009dd";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"ffed09dd";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"0c038104";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"ffc209dd";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"005109dd";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"04061810";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"0102a204";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"ffec09dd";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"96059e08";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"ac019204";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"000509dd";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"009509dd";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"fff609dd";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"560b5804";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"ffa109dd";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"9203d904";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"ffdf09dd";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"006d09dd";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"3905e11c";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"8efab308";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"f1001104";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"009d0a61";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"ffab0a61";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"20083308";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"010b8604";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"ff680a61";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"fff00a61";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"13090e08";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"a2001d04";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"fff00a61";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"ff990a61";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"00580a61";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"20030508";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"0c02f104";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"ff760a61";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"00010a61";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"5003b208";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"2800b704";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"00160a61";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"ff880a61";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"02073410";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"0902ed08";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"80045704";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"00890a61";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"ffe70a61";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"0401bd04";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"00380a61";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"ffa90a61";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"af01c504";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"ffa90a61";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"ffed0a61";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"4c016330";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"04032018";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"50022e04";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"ffa10add";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"47035c08";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"0f009a04";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"00440add";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"ffae0add";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"31016c04";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"fff60add";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"bf012804";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"00190add";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"00930add";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"82036608";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"560c8e04";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"ff7b0add";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"00230add";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"3a009508";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"0702c204";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"00070add";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"00760add";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"1407b104";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"ff8f0add";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"00300add";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"8efab304";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"00280add";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"140af708";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"b90cd804";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"ff690add";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"ffd90add";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"00030add";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"3905e114";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"8efab304";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"00250b69";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"0109e408";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"200ab604";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"ff690b69";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"fffc0b69";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"ae008d04";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"00470b69";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"ffc10b69";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"1603c614";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"0f04c40c";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"4702f504";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"ffb50b69";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"c3006c04";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"00750b69";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"00000b69";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"7a06ce04";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"ff810b69";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"00140b69";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"04048710";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"01036504";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"fffa0b69";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"cc06de08";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"8300fe04";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"00290b69";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"00900b69";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"001b0b69";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"2b01b708";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"2205e904";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"fffe0b69";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"00640b69";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"f6037604";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"ffa10b69";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"ffee0b69";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"50052118";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"63000108";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"8efd0404";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"00730be1";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"ffc80be1";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"660e9b0c";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"1407b108";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"21002104";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"ffca0be1";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"ff6b0be1";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"ffe10be1";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"00270be1";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"2005630c";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"1804c508";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"e504ec04";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"ff850be1";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"ffe80be1";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"001b0be1";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"0103b008";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"5c04ae04";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"ff9e0be1";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"00050be1";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"100bb00c";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"4f05bc08";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"09033704";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"00890be1";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"00040be1";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"fff20be1";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"ffcd0be1";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"ee03e60c";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"b0004304";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"00370c55";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"5006f804";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"ff6c0c55";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"ffe00c55";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"04030118";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"0205ef10";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"2003af04";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"fff30c55";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"e500cd04";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"00170c55";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"2c034504";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"00880c55";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"002a0c55";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"30003204";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"000e0c55";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"ffbd0c55";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"c604c80c";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"6400d508";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"6d03ad04";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"00640c55";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"000c0c55";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"ffc00c55";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"3f0f0708";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"9204b704";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"ff800c55";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"fff70c55";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"00130c55";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"4c016328";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"9f02a01c";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"0105230c";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"a4089f08";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"07037604";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"ffa80cb9";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"fff20cb9";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"00360cb9";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"5b02870c";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"4e077b08";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"82020604";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"00180cb9";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"00830cb9";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"fff90cb9";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"ffec0cb9";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"1f034008";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"a5043a04";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"ffd30cb9";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"00370cb9";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"ff960cb9";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"b0004304";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"002d0cb9";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"6a085a04";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"ff700cb9";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"ffee0cb9";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"3905e110";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"8efbd604";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"001e0d15";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"0109e408";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"ee09f004";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"ff700d15";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"ffd80d15";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"00000d15";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"04032010";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"56013a04";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"ffe00d15";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"1402c204";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"00050d15";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"0c00d204";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"001b0d15";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"007a0d15";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"82040c08";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"02022704";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"ffec0d15";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"ff8f0d15";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"33018f04";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"00500d15";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"ffda0d15";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"2005a118";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"19015710";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"0f02eb08";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"8c00c604";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"00600d71";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"ffe90d71";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"a1017104";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"ffec0d71";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"ff990d71";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"6008ad04";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"ff740d71";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"ffeb0d71";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"5b00aa0c";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"3f069c04";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"fff70d71";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"0404dc04";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"00780d71";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"00240d71";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"6a076b04";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"ffa50d71";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"05025f04";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"004e0d71";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"ffdc0d71";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"4705c018";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"19016c10";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"03009608";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"d2009c04";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"005d0dc5";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"00070dc5";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"9107e804";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"ff940dc5";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"000e0dc5";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"3c080c04";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"ff770dc5";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"ffee0dc5";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"5b00ee0c";
		wait for Clk_period;
		Addr <=  "0001101101001";
		Trees_din <= x"3f081804";
		wait for Clk_period;
		Addr <=  "0001101101010";
		Trees_din <= x"00060dc5";
		wait for Clk_period;
		Addr <=  "0001101101011";
		Trees_din <= x"12055f04";
		wait for Clk_period;
		Addr <=  "0001101101100";
		Trees_din <= x"00720dc5";
		wait for Clk_period;
		Addr <=  "0001101101101";
		Trees_din <= x"001f0dc5";
		wait for Clk_period;
		Addr <=  "0001101101110";
		Trees_din <= x"010a3904";
		wait for Clk_period;
		Addr <=  "0001101101111";
		Trees_din <= x"ffba0dc5";
		wait for Clk_period;
		Addr <=  "0001101110000";
		Trees_din <= x"00170dc5";
		wait for Clk_period;
		Addr <=  "0001101110001";
		Trees_din <= x"20057910";
		wait for Clk_period;
		Addr <=  "0001101110010";
		Trees_din <= x"63000104";
		wait for Clk_period;
		Addr <=  "0001101110011";
		Trees_din <= x"00210e09";
		wait for Clk_period;
		Addr <=  "0001101110100";
		Trees_din <= x"4c009208";
		wait for Clk_period;
		Addr <=  "0001101110101";
		Trees_din <= x"4e03f204";
		wait for Clk_period;
		Addr <=  "0001101110110";
		Trees_din <= x"00280e09";
		wait for Clk_period;
		Addr <=  "0001101110111";
		Trees_din <= x"ffc00e09";
		wait for Clk_period;
		Addr <=  "0001101111000";
		Trees_din <= x"ff800e09";
		wait for Clk_period;
		Addr <=  "0001101111001";
		Trees_din <= x"7c068308";
		wait for Clk_period;
		Addr <=  "0001101111010";
		Trees_din <= x"3c062e04";
		wait for Clk_period;
		Addr <=  "0001101111011";
		Trees_din <= x"ffab0e09";
		wait for Clk_period;
		Addr <=  "0001101111100";
		Trees_din <= x"001a0e09";
		wait for Clk_period;
		Addr <=  "0001101111101";
		Trees_din <= x"1d06d008";
		wait for Clk_period;
		Addr <=  "0001101111110";
		Trees_din <= x"0b0b1904";
		wait for Clk_period;
		Addr <=  "0001101111111";
		Trees_din <= x"006e0e09";
		wait for Clk_period;
		Addr <=  "0001110000000";
		Trees_din <= x"000d0e09";
		wait for Clk_period;
		Addr <=  "0001110000001";
		Trees_din <= x"fff00e09";
		wait for Clk_period;
		Addr <=  "0001110000010";
		Trees_din <= x"3c057b0c";
		wait for Clk_period;
		Addr <=  "0001110000011";
		Trees_din <= x"a4089f08";
		wait for Clk_period;
		Addr <=  "0001110000100";
		Trees_din <= x"fe000b04";
		wait for Clk_period;
		Addr <=  "0001110000101";
		Trees_din <= x"fff30e4d";
		wait for Clk_period;
		Addr <=  "0001110000110";
		Trees_din <= x"ff830e4d";
		wait for Clk_period;
		Addr <=  "0001110000111";
		Trees_din <= x"00140e4d";
		wait for Clk_period;
		Addr <=  "0001110001000";
		Trees_din <= x"3302950c";
		wait for Clk_period;
		Addr <=  "0001110001001";
		Trees_din <= x"04028304";
		wait for Clk_period;
		Addr <=  "0001110001010";
		Trees_din <= x"006f0e4d";
		wait for Clk_period;
		Addr <=  "0001110001011";
		Trees_din <= x"14065a04";
		wait for Clk_period;
		Addr <=  "0001110001100";
		Trees_din <= x"ffea0e4d";
		wait for Clk_period;
		Addr <=  "0001110001101";
		Trees_din <= x"00410e4d";
		wait for Clk_period;
		Addr <=  "0001110001110";
		Trees_din <= x"7a067308";
		wait for Clk_period;
		Addr <=  "0001110001111";
		Trees_din <= x"3e034a04";
		wait for Clk_period;
		Addr <=  "0001110010000";
		Trees_din <= x"ffa90e4d";
		wait for Clk_period;
		Addr <=  "0001110010001";
		Trees_din <= x"fff10e4d";
		wait for Clk_period;
		Addr <=  "0001110010010";
		Trees_din <= x"00190e4d";
		wait for Clk_period;
		Addr <=  "0001110010011";
		Trees_din <= x"4705c014";
		wait for Clk_period;
		Addr <=  "0001110010100";
		Trees_din <= x"a504a908";
		wait for Clk_period;
		Addr <=  "0001110010101";
		Trees_din <= x"3f080004";
		wait for Clk_period;
		Addr <=  "0001110010110";
		Trees_din <= x"ff840e91";
		wait for Clk_period;
		Addr <=  "0001110010111";
		Trees_din <= x"ffe70e91";
		wait for Clk_period;
		Addr <=  "0001110011000";
		Trees_din <= x"19016c08";
		wait for Clk_period;
		Addr <=  "0001110011001";
		Trees_din <= x"7400ef04";
		wait for Clk_period;
		Addr <=  "0001110011010";
		Trees_din <= x"00470e91";
		wait for Clk_period;
		Addr <=  "0001110011011";
		Trees_din <= x"fffe0e91";
		wait for Clk_period;
		Addr <=  "0001110011100";
		Trees_din <= x"ffb90e91";
		wait for Clk_period;
		Addr <=  "0001110011101";
		Trees_din <= x"5b009808";
		wait for Clk_period;
		Addr <=  "0001110011110";
		Trees_din <= x"07038404";
		wait for Clk_period;
		Addr <=  "0001110011111";
		Trees_din <= x"00140e91";
		wait for Clk_period;
		Addr <=  "0001110100000";
		Trees_din <= x"00660e91";
		wait for Clk_period;
		Addr <=  "0001110100001";
		Trees_din <= x"6a076b04";
		wait for Clk_period;
		Addr <=  "0001110100010";
		Trees_din <= x"ffc60e91";
		wait for Clk_period;
		Addr <=  "0001110100011";
		Trees_din <= x"00180e91";
		wait for Clk_period;
		Addr <=  "0001110100100";
		Trees_din <= x"2004f10c";
		wait for Clk_period;
		Addr <=  "0001110100101";
		Trees_din <= x"8efde604";
		wait for Clk_period;
		Addr <=  "0001110100110";
		Trees_din <= x"00100ec5";
		wait for Clk_period;
		Addr <=  "0001110100111";
		Trees_din <= x"b909e704";
		wait for Clk_period;
		Addr <=  "0001110101000";
		Trees_din <= x"ff860ec5";
		wait for Clk_period;
		Addr <=  "0001110101001";
		Trees_din <= x"ffe50ec5";
		wait for Clk_period;
		Addr <=  "0001110101010";
		Trees_din <= x"0103b804";
		wait for Clk_period;
		Addr <=  "0001110101011";
		Trees_din <= x"ffbc0ec5";
		wait for Clk_period;
		Addr <=  "0001110101100";
		Trees_din <= x"d4045704";
		wait for Clk_period;
		Addr <=  "0001110101101";
		Trees_din <= x"ffee0ec5";
		wait for Clk_period;
		Addr <=  "0001110101110";
		Trees_din <= x"ae031604";
		wait for Clk_period;
		Addr <=  "0001110101111";
		Trees_din <= x"00620ec5";
		wait for Clk_period;
		Addr <=  "0001110110000";
		Trees_din <= x"00010ec5";
		wait for Clk_period;
		Addr <=  "0001110110001";
		Trees_din <= x"3c062e0c";
		wait for Clk_period;
		Addr <=  "0001110110010";
		Trees_din <= x"a4089f08";
		wait for Clk_period;
		Addr <=  "0001110110011";
		Trees_din <= x"7700b204";
		wait for Clk_period;
		Addr <=  "0001110110100";
		Trees_din <= x"ffe80ef9";
		wait for Clk_period;
		Addr <=  "0001110110101";
		Trees_din <= x"ff8e0ef9";
		wait for Clk_period;
		Addr <=  "0001110110110";
		Trees_din <= x"00140ef9";
		wait for Clk_period;
		Addr <=  "0001110110111";
		Trees_din <= x"33029508";
		wait for Clk_period;
		Addr <=  "0001110111000";
		Trees_din <= x"2b01ab04";
		wait for Clk_period;
		Addr <=  "0001110111001";
		Trees_din <= x"005f0ef9";
		wait for Clk_period;
		Addr <=  "0001110111010";
		Trees_din <= x"00160ef9";
		wait for Clk_period;
		Addr <=  "0001110111011";
		Trees_din <= x"50090204";
		wait for Clk_period;
		Addr <=  "0001110111100";
		Trees_din <= x"ffb60ef9";
		wait for Clk_period;
		Addr <=  "0001110111101";
		Trees_din <= x"00100ef9";
		wait for Clk_period;
		Addr <=  "0001110111110";
		Trees_din <= x"3f0bf914";
		wait for Clk_period;
		Addr <=  "0001110111111";
		Trees_din <= x"1305c408";
		wait for Clk_period;
		Addr <=  "0001111000000";
		Trees_din <= x"7400fd04";
		wait for Clk_period;
		Addr <=  "0001111000001";
		Trees_din <= x"ffef0f2d";
		wait for Clk_period;
		Addr <=  "0001111000010";
		Trees_din <= x"ff920f2d";
		wait for Clk_period;
		Addr <=  "0001111000011";
		Trees_din <= x"6c040d08";
		wait for Clk_period;
		Addr <=  "0001111000100";
		Trees_din <= x"3c051c04";
		wait for Clk_period;
		Addr <=  "0001111000101";
		Trees_din <= x"00020f2d";
		wait for Clk_period;
		Addr <=  "0001111000110";
		Trees_din <= x"00430f2d";
		wait for Clk_period;
		Addr <=  "0001111000111";
		Trees_din <= x"ffce0f2d";
		wait for Clk_period;
		Addr <=  "0001111001000";
		Trees_din <= x"8b03c704";
		wait for Clk_period;
		Addr <=  "0001111001001";
		Trees_din <= x"00030f2d";
		wait for Clk_period;
		Addr <=  "0001111001010";
		Trees_din <= x"00520f2d";
		wait for Clk_period;
		Addr <=  "0001111001011";
		Trees_din <= x"3905e108";
		wait for Clk_period;
		Addr <=  "0001111001100";
		Trees_din <= x"3106c304";
		wait for Clk_period;
		Addr <=  "0001111001101";
		Trees_din <= x"ff9a0f61";
		wait for Clk_period;
		Addr <=  "0001111001110";
		Trees_din <= x"ffff0f61";
		wait for Clk_period;
		Addr <=  "0001111001111";
		Trees_din <= x"1603c608";
		wait for Clk_period;
		Addr <=  "0001111010000";
		Trees_din <= x"0f04c404";
		wait for Clk_period;
		Addr <=  "0001111010001";
		Trees_din <= x"00130f61";
		wait for Clk_period;
		Addr <=  "0001111010010";
		Trees_din <= x"ffc50f61";
		wait for Clk_period;
		Addr <=  "0001111010011";
		Trees_din <= x"04048708";
		wait for Clk_period;
		Addr <=  "0001111010100";
		Trees_din <= x"02025f04";
		wait for Clk_period;
		Addr <=  "0001111010101";
		Trees_din <= x"005f0f61";
		wait for Clk_period;
		Addr <=  "0001111010110";
		Trees_din <= x"00130f61";
		wait for Clk_period;
		Addr <=  "0001111010111";
		Trees_din <= x"fff90f61";
		wait for Clk_period;
		Addr <=  "0001111011000";
		Trees_din <= x"20057908";
		wait for Clk_period;
		Addr <=  "0001111011001";
		Trees_din <= x"a504a904";
		wait for Clk_period;
		Addr <=  "0001111011010";
		Trees_din <= x"ffa40f85";
		wait for Clk_period;
		Addr <=  "0001111011011";
		Trees_din <= x"fffc0f85";
		wait for Clk_period;
		Addr <=  "0001111011100";
		Trees_din <= x"7c068304";
		wait for Clk_period;
		Addr <=  "0001111011101";
		Trees_din <= x"ffde0f85";
		wait for Clk_period;
		Addr <=  "0001111011110";
		Trees_din <= x"01081b04";
		wait for Clk_period;
		Addr <=  "0001111011111";
		Trees_din <= x"00010f85";
		wait for Clk_period;
		Addr <=  "0001111100000";
		Trees_din <= x"004d0f85";
		wait for Clk_period;
		Addr <=  "0001111100001";
		Trees_din <= x"3c062e0c";
		wait for Clk_period;
		Addr <=  "0001111100010";
		Trees_din <= x"7700b208";
		wait for Clk_period;
		Addr <=  "0001111100011";
		Trees_din <= x"9a022a04";
		wait for Clk_period;
		Addr <=  "0001111100100";
		Trees_din <= x"ffeb0fb1";
		wait for Clk_period;
		Addr <=  "0001111100101";
		Trees_din <= x"00180fb1";
		wait for Clk_period;
		Addr <=  "0001111100110";
		Trees_din <= x"ffa90fb1";
		wait for Clk_period;
		Addr <=  "0001111100111";
		Trees_din <= x"4e062008";
		wait for Clk_period;
		Addr <=  "0001111101000";
		Trees_din <= x"3301ff04";
		wait for Clk_period;
		Addr <=  "0001111101001";
		Trees_din <= x"00570fb1";
		wait for Clk_period;
		Addr <=  "0001111101010";
		Trees_din <= x"00060fb1";
		wait for Clk_period;
		Addr <=  "0001111101011";
		Trees_din <= x"ffd90fb1";
		wait for Clk_period;
		Addr <=  "0001111101100";
		Trees_din <= x"14065a0c";
		wait for Clk_period;
		Addr <=  "0001111101101";
		Trees_din <= x"8b07ea08";
		wait for Clk_period;
		Addr <=  "0001111101110";
		Trees_din <= x"9a03c204";
		wait for Clk_period;
		Addr <=  "0001111101111";
		Trees_din <= x"ffa60fd5";
		wait for Clk_period;
		Addr <=  "0001111110000";
		Trees_din <= x"fff70fd5";
		wait for Clk_period;
		Addr <=  "0001111110001";
		Trees_din <= x"00220fd5";
		wait for Clk_period;
		Addr <=  "0001111110010";
		Trees_din <= x"0d041204";
		wait for Clk_period;
		Addr <=  "0001111110011";
		Trees_din <= x"00010fd5";
		wait for Clk_period;
		Addr <=  "0001111110100";
		Trees_din <= x"00470fd5";
		wait for Clk_period;
		Addr <=  "0001111110101";
		Trees_din <= x"3f0f0710";
		wait for Clk_period;
		Addr <=  "0001111110110";
		Trees_din <= x"3302190c";
		wait for Clk_period;
		Addr <=  "0001111110111";
		Trees_din <= x"3c062e08";
		wait for Clk_period;
		Addr <=  "0001111111000";
		Trees_din <= x"7700ac04";
		wait for Clk_period;
		Addr <=  "0001111111001";
		Trees_din <= x"00120ff9";
		wait for Clk_period;
		Addr <=  "0001111111010";
		Trees_din <= x"ffbd0ff9";
		wait for Clk_period;
		Addr <=  "0001111111011";
		Trees_din <= x"00370ff9";
		wait for Clk_period;
		Addr <=  "0001111111100";
		Trees_din <= x"ffb00ff9";
		wait for Clk_period;
		Addr <=  "0001111111101";
		Trees_din <= x"00420ff9";
		wait for Clk_period;
		Addr <=  "0001111111110";
		Trees_din <= x"470a450c";
		wait for Clk_period;
		Addr <=  "0001111111111";
		Trees_din <= x"c3006504";
		wait for Clk_period;
		Addr <=  "0010000000000";
		Trees_din <= x"0011101d";
		wait for Clk_period;
		Addr <=  "0010000000001";
		Trees_din <= x"0300d104";
		wait for Clk_period;
		Addr <=  "0010000000010";
		Trees_din <= x"fff5101d";
		wait for Clk_period;
		Addr <=  "0010000000011";
		Trees_din <= x"ffb1101d";
		wait for Clk_period;
		Addr <=  "0010000000100";
		Trees_din <= x"0401ea04";
		wait for Clk_period;
		Addr <=  "0010000000101";
		Trees_din <= x"0044101d";
		wait for Clk_period;
		Addr <=  "0010000000110";
		Trees_din <= x"0011101d";
		wait for Clk_period;
		Addr <=  "0010000000111";
		Trees_din <= x"ae02990c";
		wait for Clk_period;
		Addr <=  "0010000001000";
		Trees_din <= x"3d00c908";
		wait for Clk_period;
		Addr <=  "0010000001001";
		Trees_din <= x"04033a04";
		wait for Clk_period;
		Addr <=  "0010000001010";
		Trees_din <= x"004b1041";
		wait for Clk_period;
		Addr <=  "0010000001011";
		Trees_din <= x"00081041";
		wait for Clk_period;
		Addr <=  "0010000001100";
		Trees_din <= x"ffe11041";
		wait for Clk_period;
		Addr <=  "0010000001101";
		Trees_din <= x"20056304";
		wait for Clk_period;
		Addr <=  "0010000001110";
		Trees_din <= x"ffb51041";
		wait for Clk_period;
		Addr <=  "0010000001111";
		Trees_din <= x"fff51041";
		wait for Clk_period;
		Addr <=  "0010000010000";
		Trees_din <= x"39064f08";
		wait for Clk_period;
		Addr <=  "0010000010001";
		Trees_din <= x"2b01b304";
		wait for Clk_period;
		Addr <=  "0010000010010";
		Trees_din <= x"fff9105d";
		wait for Clk_period;
		Addr <=  "0010000010011";
		Trees_din <= x"ffb5105d";
		wait for Clk_period;
		Addr <=  "0010000010100";
		Trees_din <= x"05029e04";
		wait for Clk_period;
		Addr <=  "0010000010101";
		Trees_din <= x"003c105d";
		wait for Clk_period;
		Addr <=  "0010000010110";
		Trees_din <= x"fff1105d";
		wait for Clk_period;
		Addr <=  "0010000010111";
		Trees_din <= x"9f02a010";
		wait for Clk_period;
		Addr <=  "0010000011000";
		Trees_din <= x"0d043908";
		wait for Clk_period;
		Addr <=  "0010000011001";
		Trees_din <= x"8501c504";
		wait for Clk_period;
		Addr <=  "0010000011010";
		Trees_din <= x"00121081";
		wait for Clk_period;
		Addr <=  "0010000011011";
		Trees_din <= x"ffd21081";
		wait for Clk_period;
		Addr <=  "0010000011100";
		Trees_din <= x"07045d04";
		wait for Clk_period;
		Addr <=  "0010000011101";
		Trees_din <= x"00111081";
		wait for Clk_period;
		Addr <=  "0010000011110";
		Trees_din <= x"00461081";
		wait for Clk_period;
		Addr <=  "0010000011111";
		Trees_din <= x"ffc81081";
		wait for Clk_period;
		Addr <=  "0010000100000";
		Trees_din <= x"0403010c";
		wait for Clk_period;
		Addr <=  "0010000100001";
		Trees_din <= x"6a052e04";
		wait for Clk_period;
		Addr <=  "0010000100010";
		Trees_din <= x"ffee10a5";
		wait for Clk_period;
		Addr <=  "0010000100011";
		Trees_din <= x"56045304";
		wait for Clk_period;
		Addr <=  "0010000100100";
		Trees_din <= x"001110a5";
		wait for Clk_period;
		Addr <=  "0010000100101";
		Trees_din <= x"004510a5";
		wait for Clk_period;
		Addr <=  "0010000100110";
		Trees_din <= x"3e077b04";
		wait for Clk_period;
		Addr <=  "0010000100111";
		Trees_din <= x"ffbe10a5";
		wait for Clk_period;
		Addr <=  "0010000101000";
		Trees_din <= x"000410a5";
		wait for Clk_period;
		Addr <=  "0010000101001";
		Trees_din <= x"ae029908";
		wait for Clk_period;
		Addr <=  "0010000101010";
		Trees_din <= x"3c057b04";
		wait for Clk_period;
		Addr <=  "0010000101011";
		Trees_din <= x"ffed10b9";
		wait for Clk_period;
		Addr <=  "0010000101100";
		Trees_din <= x"003810b9";
		wait for Clk_period;
		Addr <=  "0010000101101";
		Trees_din <= x"ffce10b9";
		wait for Clk_period;
		Addr <=  "0010000101110";
		Trees_din <= x"04030108";
		wait for Clk_period;
		Addr <=  "0010000101111";
		Trees_din <= x"30015704";
		wait for Clk_period;
		Addr <=  "0010000110000";
		Trees_din <= x"003610d5";
		wait for Clk_period;
		Addr <=  "0010000110001";
		Trees_din <= x"ffef10d5";
		wait for Clk_period;
		Addr <=  "0010000110010";
		Trees_din <= x"3e077b04";
		wait for Clk_period;
		Addr <=  "0010000110011";
		Trees_din <= x"ffc410d5";
		wait for Clk_period;
		Addr <=  "0010000110100";
		Trees_din <= x"000110d5";
		wait for Clk_period;
		Addr <=  "0010000110101";
		Trees_din <= x"0109120c";
		wait for Clk_period;
		Addr <=  "0010000110110";
		Trees_din <= x"7400ef04";
		wait for Clk_period;
		Addr <=  "0010000110111";
		Trees_din <= x"000c10f9";
		wait for Clk_period;
		Addr <=  "0010000111000";
		Trees_din <= x"13042a04";
		wait for Clk_period;
		Addr <=  "0010000111001";
		Trees_din <= x"ffc010f9";
		wait for Clk_period;
		Addr <=  "0010000111010";
		Trees_din <= x"fff210f9";
		wait for Clk_period;
		Addr <=  "0010000111011";
		Trees_din <= x"40017b04";
		wait for Clk_period;
		Addr <=  "0010000111100";
		Trees_din <= x"000610f9";
		wait for Clk_period;
		Addr <=  "0010000111101";
		Trees_din <= x"003710f9";
		wait for Clk_period;
		Addr <=  "0010000111110";
		Trees_din <= x"3f0f0708";
		wait for Clk_period;
		Addr <=  "0010000111111";
		Trees_din <= x"1305c404";
		wait for Clk_period;
		Addr <=  "0010001000000";
		Trees_din <= x"ffc8110d";
		wait for Clk_period;
		Addr <=  "0010001000001";
		Trees_din <= x"000e110d";
		wait for Clk_period;
		Addr <=  "0010001000010";
		Trees_din <= x"0033110d";
		wait for Clk_period;
		Addr <=  "0010001000011";
		Trees_din <= x"b9061a04";
		wait for Clk_period;
		Addr <=  "0010001000100";
		Trees_din <= x"ffd61121";
		wait for Clk_period;
		Addr <=  "0010001000101";
		Trees_din <= x"0d041204";
		wait for Clk_period;
		Addr <=  "0010001000110";
		Trees_din <= x"ffee1121";
		wait for Clk_period;
		Addr <=  "0010001000111";
		Trees_din <= x"00311121";
		wait for Clk_period;
		Addr <=  "0010001001000";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  4
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"1207dc4c";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"0509792c";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"420adb1c";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"180a1c10";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"08000b08";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"4d02fc04";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"ff6e0125";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"02890125";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"460a3a04";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"ff540125";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"00200125";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"30038f08";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"48039504";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"039c0125";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"00120125";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"ff5f0125";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"08019108";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"6601a204";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"00270125";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"03710125";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"0000f504";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"00270125";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"ff890125";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"b101f408";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"13070804";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"ff5c0125";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"00b20125";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"5a017b08";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"0801b304";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"013c0125";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"ff850125";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"02013a08";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"08026904";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"013c0125";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"ff9d0125";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"2f042e04";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"04090125";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"00b20125";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"03032c20";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"0507d118";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"460a1310";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"1309db08";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"b8000604";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"00e20125";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"ff640125";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"57025c04";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"ff810125";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"026a0125";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"16068f04";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"03270125";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"ff9d0125";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"0902de04";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"03ae0125";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"00270125";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"2b04d218";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"c000a308";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"2600af04";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"02360125";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"ff730125";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"7907f708";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"f2046d04";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"041d0125";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"01700125";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"0305ab04";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"ff9d0125";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"013c0125";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"0800b408";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"42036604";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"00b20125";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"03220125";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"02088304";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"ff610125";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"013c0125";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"a805b754";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"1208812c";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"130e641c";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"310c990c";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"660e9b08";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"420a6104";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"ff570289";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"001f0289";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"00af0289";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"0701ed08";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"57033a04";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"ff9a0289";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"01d30289";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"7d030a04";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"ff690289";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"00370289";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"3e05450c";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"0802a308";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"7a023f04";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"02530289";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"00ad0289";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"ffa30289";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"ff750289";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"18033b10";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"74006a08";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"0700eb04";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"012c0289";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"00190289";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"9f084f04";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"ff5b0289";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"002f0289";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"65003c08";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"53020304";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"003a0289";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"ff790289";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"7604a408";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"2905fe04";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"01cd0289";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"00180289";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"06015b04";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"00ff0289";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"ff7c0289";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"0203b138";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"0504c41c";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"0f0c8610";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"2e079a08";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"ad0bad04";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"ff580289";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"003b0289";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"0f044d04";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"ff910289";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"018b0289";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"e8094704";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"01b20289";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"f0000804";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"00320289";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"ff810289";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"dc045410";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"4605f308";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"34077f04";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"ff630289";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"00ae0289";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"0f04c404";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"ff7e0289";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"01a90289";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"8207f508";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"6f02b704";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"01c90289";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"ffcb0289";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"ff730289";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"05020a10";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"08008408";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"1202c804";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"ff9f0289";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"01920289";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"98103d04";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"ff5d0289";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"00ab0289";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"0906680c";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"3e0d2d08";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"0a0b2104";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"01b60289";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"ff920289";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"ff840289";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"9808a008";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"74007004";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"009f0289";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"ff610289";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"013e0289";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"a805b750";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"1208812c";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"130cb91c";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"310b7510";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"2c004708";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"e801ce04";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"016803e5";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"ff6403e5";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"460ef104";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"ff5a03e5";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"001e03e5";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"40015908";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"b9076504";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"015803e5";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"ff8903e5";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"ff6803e5";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"3e05450c";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"b101f404";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"ff9103e5";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"05018c04";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"002903e5";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"019b03e5";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"ff6d03e5";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"18033b10";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"74006a08";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"2804dd04";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"000e03e5";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"00f903e5";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"9f084f04";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"ff6203e5";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"002a03e5";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"ee013a04";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"ff7d03e5";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"15052c08";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"48057404";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"014003e5";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"ff9e03e5";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"b0052104";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"ff9203e5";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"002103e5";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"05044438";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"0205031c";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"0f0c8610";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"2e079a08";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"d8001f04";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"001a03e5";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"ff6003e5";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"40004d04";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"014203e5";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"ff8e03e5";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"53026404";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"014503e5";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"b7107504";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"ff8103e5";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"002f03e5";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"1205770c";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"5300c708";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"0502e504";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"ffaa03e5";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"010803e5";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"ff6603e5";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"79041d08";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"0302a204";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"005003e5";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"014603e5";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"0a023c04";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"003703e5";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"ff8e03e5";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"0906421c";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"e20ae810";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"2f045608";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"48082f04";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"013a03e5";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"ff8f03e5";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"0f04c404";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"ff6f03e5";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"00e503e5";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"0c006a08";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"5a070004";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"000303e5";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"010003e5";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"ff6c03e5";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"0207b608";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"6a0a0504";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"ff5c03e5";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"00e103e5";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"010903e5";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"0b03c640";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"1208ba24";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"420a611c";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"05097910";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"7f000808";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"56013e04";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"00da0509";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"ff890509";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"740cd004";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"ff5c0509";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"ffca0509";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"9f070904";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"ff6d0509";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"7f021804";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"00e30509";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"002a0509";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"7b014d04";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"012c0509";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"ff8d0509";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"4b028708";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"87128f04";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"ff620509";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"00100509";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"7f009308";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"0903f904";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"01050509";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"00480509";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"4c01ec08";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"2b00ee04";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"00c50509";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"ffff0509";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"ff740509";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"0f03df30";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"7400c314";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"7504dc10";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"45034b08";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"4c001b04";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"006f0509";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"ff710509";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"1903d104";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"011a0509";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"fff20509";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"ff690509";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"130b7910";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"310ef308";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"0f03cd04";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"ff5b0509";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"000b0509";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"52000404";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"ffac0509";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"00910509";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"1605b508";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"b6033a04";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"01070509";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"00090509";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"ff770509";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"16077c18";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"7f039210";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"82063f08";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"93001504";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"ff850509";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"01010509";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"1207b204";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"ff6c0509";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"00b40509";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"b8000b04";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"006a0509";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"ff6e0509";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"05092408";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"2807ad04";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"ff600509";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"00710509";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"00b20509";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"0b03c644";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"1208ba28";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"420a6120";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"05089d10";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"7f000808";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"5e02d904";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"ff910645";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"00b50645";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"82001004";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"ffde0645";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"ff5f0645";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"7a00a108";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"7b014d04";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"010a0645";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"ffaa0645";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"9b013804";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"fffc0645";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"ff6e0645";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"7b014d04";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"01020645";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"ff960645";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"4b028708";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"bf0b3e04";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"ff670645";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"00090645";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"5a00fb08";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"11029004";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"fffc0645";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"ff940645";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"45032104";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"ffd00645";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"0904d504";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"00e20645";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"fff90645";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"0503c534";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"12048d1c";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"1309860c";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"f00a7808";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"50000404";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"00040645";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"ff5f0645";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"00650645";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"fd039708";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"86013004";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"01030645";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"fff40645";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"fa003904";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"002d0645";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"ff6b0645";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"2203cf10";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"f5023508";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"82059e04";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"00d10645";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"ff8d0645";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"e6008904";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"fffd0645";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"ff850645";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"120e8804";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"ff660645";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"00650645";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"0f018f0c";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"7400a408";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"03061f04";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"fffc0645";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"00a40645";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"ff6b0645";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"2b061b10";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"c000cc08";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"8c004a04";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"00830645";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"ff7a0645";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"7f03b804";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"00de0645";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"ffad0645";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"4f025d04";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"ff6c0645";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"8302aa04";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"00be0645";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"ff810645";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"0b03c640";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"1208ba24";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"420a611c";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"05089d10";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"7f000808";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"9a043e04";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"ff7c0779";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"007f0779";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"82001004";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"ffea0779";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"ff610779";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"f2018908";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"80046d04";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"ff9e0779";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"00dc0779";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"ff780779";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"7b014d04";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"00e60779";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"ff9f0779";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"4b028708";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"4a000004";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"00050779";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"ff6d0779";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"7f009308";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"15044a04";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"00c90779";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"002d0779";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"90001404";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"008c0779";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"5505d504";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"ff830779";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"ffef0779";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"0f03df2c";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"7400c314";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"7504dc10";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"45034b08";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"bd05a604";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"ff7a0779";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"00410779";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"5302de04";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"00de0779";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"00100779";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"ff740779";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"130b790c";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"310ef308";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"d8000704";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"fff10779";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"ff600779";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"00250779";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"1605b508";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"b3015604";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"00bc0779";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"00090779";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"ff840779";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"1607101c";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"49058f0c";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"eb011204";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"ff8d0779";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"500cb304";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"00c60779";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"ffe30779";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"7f004f08";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"e4014e04";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"00a80779";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"ffff0779";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"c80a9604";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"ff6d0779";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"fff60779";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"0204ea08";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"cd019804";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"ffef0779";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"ff680779";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"4001cf08";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"42038504";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"00220779";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"00a90779";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"ffa20779";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"0b03c640";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"1208ba28";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"420a6120";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"05078e10";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"7f000808";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"9a043e04";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"ff8208b5";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"006a08b5";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"08003e04";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"ffd408b5";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"ff6208b5";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"7a00a108";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"80069604";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"ffca08b5";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"00db08b5";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"18066e04";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"ff7308b5";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"ffec08b5";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"7b014d04";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"00d208b5";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"ffa808b5";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"4b028708";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"1705f204";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"ff7208b5";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"fffe08b5";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"5a01ba08";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"2b005c04";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"007108b5";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"ff8a08b5";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"3402da04";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"001908b5";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"00b608b5";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"2c01712c";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"16077c20";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"79066d10";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"30038f08";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"83100c04";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"00b908b5";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"ffb708b5";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"a302db04";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"009808b5";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"ff7908b5";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"5302ff08";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"df040d04";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"ffd908b5";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"00b208b5";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"03092604";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"ff6d08b5";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"004708b5";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"94031304";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"007308b5";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"0b143d04";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"ff6a08b5";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"001208b5";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"5704ef1c";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"05060b0c";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"63002804";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"003408b5";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"27003104";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"ffe908b5";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"ff6108b5";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"2e082f08";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"42080304";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"ff6d08b5";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"006908b5";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"23040c04";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"fff408b5";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"00a108b5";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"30034d10";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"40018108";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"6a026b04";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"ffeb08b5";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"00c308b5";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"46073104";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"ff9108b5";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"005708b5";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"a0048004";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"ff7c08b5";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"ffe908b5";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"b1018e1c";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"2c007c0c";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"1e03f008";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"77012d04";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"00ca09bd";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"002009bd";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"ff7b09bd";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"420a610c";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"74007008";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"3d009704";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"00da09bd";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"ff7b09bd";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"ff6309bd";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"007209bd";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"05036330";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"e2030818";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"0702c210";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"4903fb08";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"b2037304";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"00a009bd";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"ffb609bd";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"83000404";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"ffe109bd";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"ff8409bd";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"85006704";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"003209bd";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"ff6d09bd";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"0f0c2c10";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"020acf08";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"970baf04";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"ff6609bd";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"ffe209bd";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"21013904";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"006009bd";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"ffd109bd";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"2b036f04";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"008d09bd";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"ff9c09bd";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"2b04e420";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"03013c10";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"56039508";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"1f056504";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"ffcf09bd";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"008109bd";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"7b001004";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"003e09bd";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"ff7609bd";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"a3046408";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"0a0ac004";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"00ae09bd";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"ffa609bd";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"6f024004";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"006e09bd";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"ff7909bd";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"05097910";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"2c001c08";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"72006804";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"001309bd";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"006809bd";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"97071c04";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"ff6809bd";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"001509bd";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"4f01a704";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"ffab09bd";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"009509bd";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"0b03c640";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"4100cc20";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"4203ec08";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"66057d04";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"ff720ae9";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"00170ae9";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"0d04460c";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"02054d04";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"ff8e0ae9";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"de00a604";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"00700ae9";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"001b0ae9";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"3803f904";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"00030ae9";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"7701ac04";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"00da0ae9";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"003e0ae9";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"130abc14";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"af000004";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"002a0ae9";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"03097708";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"050a2904";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"ff650ae9";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"ffeb0ae9";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"2700b704";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"00630ae9";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"ffa40ae9";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"b102c304";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"ff9c0ae9";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"d2007404";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"00840ae9";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"00210ae9";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"1203ab30";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"4f05bc1c";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"ab05080c";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"a10c2008";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"bd090c04";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"ff690ae9";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"ffe20ae9";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"00220ae9";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"3a018b08";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"53038104";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"009c0ae9";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"00140ae9";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"e0066b04";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"ff840ae9";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"000d0ae9";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"d0021c0c";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"30036f08";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"8a03a904";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"00a10ae9";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"ffea0ae9";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"ffb50ae9";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"cb011d04";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"00330ae9";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"ff750ae9";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"16077c1c";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"1e07f910";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"07055c08";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"30031204";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"00a80ae9";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"001f0ae9";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"1f057c04";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"ff860ae9";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"004d0ae9";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"4604d208";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"88002104";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"fffd0ae9";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"ff820ae9";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"007a0ae9";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"05085708";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"38082904";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"ff750ae9";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"ffdc0ae9";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"00720ae9";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"2c017154";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"0302bc28";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"2e012110";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"02076508";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"8f130304";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"ff690bfd";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"ffe60bfd";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"ab067204";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"ffe40bfd";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"005a0bfd";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"0d03af08";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"59000604";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"00330bfd";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"ff780bfd";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"07017c08";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"9802bd04";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"00180bfd";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"00b80bfd";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"c6068404";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"ffa40bfd";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"00510bfd";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"09065520";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"1605b510";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"30038f08";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"7909f004";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"00a80bfd";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"ffe60bfd";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"a302db04";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"00750bfd";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"ff8d0bfd";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"42043a08";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"fe000004";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"00050bfd";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"ff880bfd";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"28021b04";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"fffa0bfd";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"00820bfd";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"aa04ba08";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"6c036d04";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"ffce0bfd";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"00770bfd";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"ff800bfd";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"02078a24";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"2200580c";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"dc03cf04";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"ff9b0bfd";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"5703cf04";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"00170bfd";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"00a20bfd";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"5800160c";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"5301fa08";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"22018c04";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"007a0bfd";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"00020bfd";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"ff8a0bfd";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"0f0b8308";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"0b0f9104";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"ff650bfd";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"ffd90bfd";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"00090bfd";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"5802a70c";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"dc015004";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"ffcc0bfd";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"12030004";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"000d0bfd";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"00990bfd";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"ce047a04";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"ff8e0bfd";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"ffe90bfd";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"2c017160";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"0302bc30";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"18045220";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"2e033f10";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"9b07a408";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"8f130304";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"ff6b0d21";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"ffe30d21";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"c3011404";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"002e0d21";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"ff9f0d21";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"86008a08";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"3a007204";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"007e0d21";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"00210d21";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"2d00e904";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"ffea0d21";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"ffae0d21";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"d604d60c";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"50073908";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"56046d04";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"00a70d21";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"001b0d21";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"ffbf0d21";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"ff9d0d21";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"1904d71c";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"0802d30c";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"730a5008";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"a8024004";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"fff30d21";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"00a20d21";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"ffe20d21";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"0f073b08";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"4f058d04";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"ff930d21";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"003f0d21";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"7903e404";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"008d0d21";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"ffe00d21";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"8401910c";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"b1017f04";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"ffb10d21";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"8200c604";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"008f0d21";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"00240d21";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"7800f204";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"001a0d21";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"ff7e0d21";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"1f06af18";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"6f000808";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"50033d04";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"00600d21";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"ffde0d21";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"a10cc10c";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"77000f04";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"ffdd0d21";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"02091104";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"ff650d21";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"ffc70d21";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"00020d21";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"3104c30c";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"55087c08";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"56007504";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"fff60d21";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"ff730d21";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"00540d21";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"0903f10c";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"84061208";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"15025404";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"00ab0d21";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"00230d21";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"000a0d21";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"ffa80d21";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"2c010e44";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"03028b20";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"2e013a0c";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"05069404";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"ff720e0d";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"02040904";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"ffb80e0d";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"00400e0d";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"5c02460c";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"0d02a204";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"ffbb0e0d";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"5d035f04";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"00180e0d";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"009b0e0d";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"19012604";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"00050e0d";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"ffa10e0d";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"09065518";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"16068f10";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"79090f08";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"07052704";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"009e0e0d";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"00190e0d";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"0d03c404";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"ffaa0e0d";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"00350e0d";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"42056804";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"ffad0e0d";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"00550e0d";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"aa04ba08";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"6c062804";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"00080e0d";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"005b0e0d";
		wait for Clk_period;
		Addr <=  "0001101101001";
		Trees_din <= x"ff910e0d";
		wait for Clk_period;
		Addr <=  "0001101101010";
		Trees_din <= x"1f067918";
		wait for Clk_period;
		Addr <=  "0001101101011";
		Trees_din <= x"6f000808";
		wait for Clk_period;
		Addr <=  "0001101101100";
		Trees_din <= x"e4010704";
		wait for Clk_period;
		Addr <=  "0001101101101";
		Trees_din <= x"00620e0d";
		wait for Clk_period;
		Addr <=  "0001101101110";
		Trees_din <= x"ffe40e0d";
		wait for Clk_period;
		Addr <=  "0001101101111";
		Trees_din <= x"4609bd08";
		wait for Clk_period;
		Addr <=  "0001101110000";
		Trees_din <= x"ad0a7104";
		wait for Clk_period;
		Addr <=  "0001101110001";
		Trees_din <= x"ff670e0d";
		wait for Clk_period;
		Addr <=  "0001101110010";
		Trees_din <= x"fff30e0d";
		wait for Clk_period;
		Addr <=  "0001101110011";
		Trees_din <= x"4f046c04";
		wait for Clk_period;
		Addr <=  "0001101110100";
		Trees_din <= x"ffa10e0d";
		wait for Clk_period;
		Addr <=  "0001101110101";
		Trees_din <= x"004e0e0d";
		wait for Clk_period;
		Addr <=  "0001101110110";
		Trees_din <= x"0203d80c";
		wait for Clk_period;
		Addr <=  "0001101110111";
		Trees_din <= x"08006304";
		wait for Clk_period;
		Addr <=  "0001101111000";
		Trees_din <= x"00500e0d";
		wait for Clk_period;
		Addr <=  "0001101111001";
		Trees_din <= x"18052004";
		wait for Clk_period;
		Addr <=  "0001101111010";
		Trees_din <= x"ff730e0d";
		wait for Clk_period;
		Addr <=  "0001101111011";
		Trees_din <= x"001a0e0d";
		wait for Clk_period;
		Addr <=  "0001101111100";
		Trees_din <= x"0d049008";
		wait for Clk_period;
		Addr <=  "0001101111101";
		Trees_din <= x"a807c504";
		wait for Clk_period;
		Addr <=  "0001101111110";
		Trees_din <= x"ffa90e0d";
		wait for Clk_period;
		Addr <=  "0001101111111";
		Trees_din <= x"00530e0d";
		wait for Clk_period;
		Addr <=  "0001110000000";
		Trees_din <= x"86027004";
		wait for Clk_period;
		Addr <=  "0001110000001";
		Trees_din <= x"009a0e0d";
		wait for Clk_period;
		Addr <=  "0001110000010";
		Trees_din <= x"001f0e0d";
		wait for Clk_period;
		Addr <=  "0001110000011";
		Trees_din <= x"2c017150";
		wait for Clk_period;
		Addr <=  "0001110000100";
		Trees_din <= x"0302bc24";
		wait for Clk_period;
		Addr <=  "0001110000101";
		Trees_din <= x"0800710c";
		wait for Clk_period;
		Addr <=  "0001110000110";
		Trees_din <= x"7605b608";
		wait for Clk_period;
		Addr <=  "0001110000111";
		Trees_din <= x"4e03b504";
		wait for Clk_period;
		Addr <=  "0001110001000";
		Trees_din <= x"000a0ef1";
		wait for Clk_period;
		Addr <=  "0001110001001";
		Trees_din <= x"009f0ef1";
		wait for Clk_period;
		Addr <=  "0001110001010";
		Trees_din <= x"ffc20ef1";
		wait for Clk_period;
		Addr <=  "0001110001011";
		Trees_din <= x"1804520c";
		wait for Clk_period;
		Addr <=  "0001110001100";
		Trees_din <= x"42077708";
		wait for Clk_period;
		Addr <=  "0001110001101";
		Trees_din <= x"8b002204";
		wait for Clk_period;
		Addr <=  "0001110001110";
		Trees_din <= x"ffd60ef1";
		wait for Clk_period;
		Addr <=  "0001110001111";
		Trees_din <= x"ff700ef1";
		wait for Clk_period;
		Addr <=  "0001110010000";
		Trees_din <= x"00040ef1";
		wait for Clk_period;
		Addr <=  "0001110010001";
		Trees_din <= x"9f030904";
		wait for Clk_period;
		Addr <=  "0001110010010";
		Trees_din <= x"ff9c0ef1";
		wait for Clk_period;
		Addr <=  "0001110010011";
		Trees_din <= x"3501f004";
		wait for Clk_period;
		Addr <=  "0001110010100";
		Trees_din <= x"00770ef1";
		wait for Clk_period;
		Addr <=  "0001110010101";
		Trees_din <= x"ffda0ef1";
		wait for Clk_period;
		Addr <=  "0001110010110";
		Trees_din <= x"1904d71c";
		wait for Clk_period;
		Addr <=  "0001110010111";
		Trees_din <= x"0802d30c";
		wait for Clk_period;
		Addr <=  "0001110011000";
		Trees_din <= x"730a5008";
		wait for Clk_period;
		Addr <=  "0001110011001";
		Trees_din <= x"ca000f04";
		wait for Clk_period;
		Addr <=  "0001110011010";
		Trees_din <= x"00020ef1";
		wait for Clk_period;
		Addr <=  "0001110011011";
		Trees_din <= x"00990ef1";
		wait for Clk_period;
		Addr <=  "0001110011100";
		Trees_din <= x"ffea0ef1";
		wait for Clk_period;
		Addr <=  "0001110011101";
		Trees_din <= x"0f073b08";
		wait for Clk_period;
		Addr <=  "0001110011110";
		Trees_din <= x"8c006f04";
		wait for Clk_period;
		Addr <=  "0001110011111";
		Trees_din <= x"00230ef1";
		wait for Clk_period;
		Addr <=  "0001110100000";
		Trees_din <= x"ff9b0ef1";
		wait for Clk_period;
		Addr <=  "0001110100001";
		Trees_din <= x"15025404";
		wait for Clk_period;
		Addr <=  "0001110100010";
		Trees_din <= x"007e0ef1";
		wait for Clk_period;
		Addr <=  "0001110100011";
		Trees_din <= x"fff50ef1";
		wait for Clk_period;
		Addr <=  "0001110100100";
		Trees_din <= x"e400f108";
		wait for Clk_period;
		Addr <=  "0001110100101";
		Trees_din <= x"05067704";
		wait for Clk_period;
		Addr <=  "0001110100110";
		Trees_din <= x"ffec0ef1";
		wait for Clk_period;
		Addr <=  "0001110100111";
		Trees_din <= x"00730ef1";
		wait for Clk_period;
		Addr <=  "0001110101000";
		Trees_din <= x"f8049204";
		wait for Clk_period;
		Addr <=  "0001110101001";
		Trees_din <= x"ff840ef1";
		wait for Clk_period;
		Addr <=  "0001110101010";
		Trees_din <= x"00240ef1";
		wait for Clk_period;
		Addr <=  "0001110101011";
		Trees_din <= x"1f06af10";
		wait for Clk_period;
		Addr <=  "0001110101100";
		Trees_din <= x"130e640c";
		wait for Clk_period;
		Addr <=  "0001110101101";
		Trees_din <= x"5708b708";
		wait for Clk_period;
		Addr <=  "0001110101110";
		Trees_din <= x"2f002c04";
		wait for Clk_period;
		Addr <=  "0001110101111";
		Trees_din <= x"ffdc0ef1";
		wait for Clk_period;
		Addr <=  "0001110110000";
		Trees_din <= x"ff680ef1";
		wait for Clk_period;
		Addr <=  "0001110110001";
		Trees_din <= x"00020ef1";
		wait for Clk_period;
		Addr <=  "0001110110010";
		Trees_din <= x"00470ef1";
		wait for Clk_period;
		Addr <=  "0001110110011";
		Trees_din <= x"31058a0c";
		wait for Clk_period;
		Addr <=  "0001110110100";
		Trees_din <= x"0207f608";
		wait for Clk_period;
		Addr <=  "0001110110101";
		Trees_din <= x"97075704";
		wait for Clk_period;
		Addr <=  "0001110110110";
		Trees_din <= x"ff7b0ef1";
		wait for Clk_period;
		Addr <=  "0001110110111";
		Trees_din <= x"fffd0ef1";
		wait for Clk_period;
		Addr <=  "0001110111000";
		Trees_din <= x"003c0ef1";
		wait for Clk_period;
		Addr <=  "0001110111001";
		Trees_din <= x"15025404";
		wait for Clk_period;
		Addr <=  "0001110111010";
		Trees_din <= x"00910ef1";
		wait for Clk_period;
		Addr <=  "0001110111011";
		Trees_din <= x"ffeb0ef1";
		wait for Clk_period;
		Addr <=  "0001110111100";
		Trees_din <= x"b1018e18";
		wait for Clk_period;
		Addr <=  "0001110111101";
		Trees_din <= x"0800c50c";
		wait for Clk_period;
		Addr <=  "0001110111110";
		Trees_din <= x"7701c308";
		wait for Clk_period;
		Addr <=  "0001110111111";
		Trees_din <= x"0a014804";
		wait for Clk_period;
		Addr <=  "0001111000000";
		Trees_din <= x"00910fbd";
		wait for Clk_period;
		Addr <=  "0001111000001";
		Trees_din <= x"fffb0fbd";
		wait for Clk_period;
		Addr <=  "0001111000010";
		Trees_din <= x"ff9a0fbd";
		wait for Clk_period;
		Addr <=  "0001111000011";
		Trees_din <= x"4100ad08";
		wait for Clk_period;
		Addr <=  "0001111000100";
		Trees_din <= x"2e040d04";
		wait for Clk_period;
		Addr <=  "0001111000101";
		Trees_din <= x"ffa10fbd";
		wait for Clk_period;
		Addr <=  "0001111000110";
		Trees_din <= x"003a0fbd";
		wait for Clk_period;
		Addr <=  "0001111000111";
		Trees_din <= x"ff690fbd";
		wait for Clk_period;
		Addr <=  "0001111001000";
		Trees_din <= x"4f023b1c";
		wait for Clk_period;
		Addr <=  "0001111001001";
		Trees_din <= x"e202480c";
		wait for Clk_period;
		Addr <=  "0001111001010";
		Trees_din <= x"6a04e004";
		wait for Clk_period;
		Addr <=  "0001111001011";
		Trees_din <= x"ffb10fbd";
		wait for Clk_period;
		Addr <=  "0001111001100";
		Trees_din <= x"07028d04";
		wait for Clk_period;
		Addr <=  "0001111001101";
		Trees_din <= x"00720fbd";
		wait for Clk_period;
		Addr <=  "0001111001110";
		Trees_din <= x"ffdd0fbd";
		wait for Clk_period;
		Addr <=  "0001111001111";
		Trees_din <= x"0f0c8608";
		wait for Clk_period;
		Addr <=  "0001111010000";
		Trees_din <= x"66098b04";
		wait for Clk_period;
		Addr <=  "0001111010001";
		Trees_din <= x"ff720fbd";
		wait for Clk_period;
		Addr <=  "0001111010010";
		Trees_din <= x"fff50fbd";
		wait for Clk_period;
		Addr <=  "0001111010011";
		Trees_din <= x"2b01c304";
		wait for Clk_period;
		Addr <=  "0001111010100";
		Trees_din <= x"004a0fbd";
		wait for Clk_period;
		Addr <=  "0001111010101";
		Trees_din <= x"ffd90fbd";
		wait for Clk_period;
		Addr <=  "0001111010110";
		Trees_din <= x"0503da1c";
		wait for Clk_period;
		Addr <=  "0001111010111";
		Trees_din <= x"8201e610";
		wait for Clk_period;
		Addr <=  "0001111011000";
		Trees_din <= x"5200f708";
		wait for Clk_period;
		Addr <=  "0001111011001";
		Trees_din <= x"5301fa04";
		wait for Clk_period;
		Addr <=  "0001111011010";
		Trees_din <= x"00910fbd";
		wait for Clk_period;
		Addr <=  "0001111011011";
		Trees_din <= x"001c0fbd";
		wait for Clk_period;
		Addr <=  "0001111011100";
		Trees_din <= x"3702a604";
		wait for Clk_period;
		Addr <=  "0001111011101";
		Trees_din <= x"00030fbd";
		wait for Clk_period;
		Addr <=  "0001111011110";
		Trees_din <= x"ffab0fbd";
		wait for Clk_period;
		Addr <=  "0001111011111";
		Trees_din <= x"03073908";
		wait for Clk_period;
		Addr <=  "0001111100000";
		Trees_din <= x"6c02f804";
		wait for Clk_period;
		Addr <=  "0001111100001";
		Trees_din <= x"ff8c0fbd";
		wait for Clk_period;
		Addr <=  "0001111100010";
		Trees_din <= x"ffe60fbd";
		wait for Clk_period;
		Addr <=  "0001111100011";
		Trees_din <= x"00350fbd";
		wait for Clk_period;
		Addr <=  "0001111100100";
		Trees_din <= x"2301a10c";
		wait for Clk_period;
		Addr <=  "0001111100101";
		Trees_din <= x"a301be08";
		wait for Clk_period;
		Addr <=  "0001111100110";
		Trees_din <= x"0001a904";
		wait for Clk_period;
		Addr <=  "0001111100111";
		Trees_din <= x"00680fbd";
		wait for Clk_period;
		Addr <=  "0001111101000";
		Trees_din <= x"000a0fbd";
		wait for Clk_period;
		Addr <=  "0001111101001";
		Trees_din <= x"ff9e0fbd";
		wait for Clk_period;
		Addr <=  "0001111101010";
		Trees_din <= x"82062908";
		wait for Clk_period;
		Addr <=  "0001111101011";
		Trees_din <= x"cb04d104";
		wait for Clk_period;
		Addr <=  "0001111101100";
		Trees_din <= x"00960fbd";
		wait for Clk_period;
		Addr <=  "0001111101101";
		Trees_din <= x"00030fbd";
		wait for Clk_period;
		Addr <=  "0001111101110";
		Trees_din <= x"fff00fbd";
		wait for Clk_period;
		Addr <=  "0001111101111";
		Trees_din <= x"2c010e38";
		wait for Clk_period;
		Addr <=  "0001111110000";
		Trees_din <= x"0303531c";
		wait for Clk_period;
		Addr <=  "0001111110001";
		Trees_din <= x"18046410";
		wait for Clk_period;
		Addr <=  "0001111110010";
		Trees_din <= x"2e030f08";
		wait for Clk_period;
		Addr <=  "0001111110011";
		Trees_din <= x"42065404";
		wait for Clk_period;
		Addr <=  "0001111110100";
		Trees_din <= x"ff7c1079";
		wait for Clk_period;
		Addr <=  "0001111110101";
		Trees_din <= x"ffed1079";
		wait for Clk_period;
		Addr <=  "0001111110110";
		Trees_din <= x"86008604";
		wait for Clk_period;
		Addr <=  "0001111110111";
		Trees_din <= x"004e1079";
		wait for Clk_period;
		Addr <=  "0001111111000";
		Trees_din <= x"fff01079";
		wait for Clk_period;
		Addr <=  "0001111111001";
		Trees_din <= x"d604d608";
		wait for Clk_period;
		Addr <=  "0001111111010";
		Trees_din <= x"56046d04";
		wait for Clk_period;
		Addr <=  "0001111111011";
		Trees_din <= x"00871079";
		wait for Clk_period;
		Addr <=  "0001111111100";
		Trees_din <= x"00011079";
		wait for Clk_period;
		Addr <=  "0001111111101";
		Trees_din <= x"ffcc1079";
		wait for Clk_period;
		Addr <=  "0001111111110";
		Trees_din <= x"1904d710";
		wait for Clk_period;
		Addr <=  "0001111111111";
		Trees_din <= x"0705270c";
		wait for Clk_period;
		Addr <=  "0010000000000";
		Trees_din <= x"1e086208";
		wait for Clk_period;
		Addr <=  "0010000000001";
		Trees_din <= x"1201fd04";
		wait for Clk_period;
		Addr <=  "0010000000010";
		Trees_din <= x"001b1079";
		wait for Clk_period;
		Addr <=  "0010000000011";
		Trees_din <= x"00961079";
		wait for Clk_period;
		Addr <=  "0010000000100";
		Trees_din <= x"fff51079";
		wait for Clk_period;
		Addr <=  "0010000000101";
		Trees_din <= x"fffd1079";
		wait for Clk_period;
		Addr <=  "0010000000110";
		Trees_din <= x"84019104";
		wait for Clk_period;
		Addr <=  "0010000000111";
		Trees_din <= x"004c1079";
		wait for Clk_period;
		Addr <=  "0010000001000";
		Trees_din <= x"8f045d04";
		wait for Clk_period;
		Addr <=  "0010000001001";
		Trees_din <= x"ffa01079";
		wait for Clk_period;
		Addr <=  "0010000001010";
		Trees_din <= x"fff31079";
		wait for Clk_period;
		Addr <=  "0010000001011";
		Trees_din <= x"1f067910";
		wait for Clk_period;
		Addr <=  "0010000001100";
		Trees_din <= x"6f000804";
		wait for Clk_period;
		Addr <=  "0010000001101";
		Trees_din <= x"002f1079";
		wait for Clk_period;
		Addr <=  "0010000001110";
		Trees_din <= x"130cb908";
		wait for Clk_period;
		Addr <=  "0010000001111";
		Trees_din <= x"02095a04";
		wait for Clk_period;
		Addr <=  "0010000010000";
		Trees_din <= x"ff6c1079";
		wait for Clk_period;
		Addr <=  "0010000010001";
		Trees_din <= x"ffeb1079";
		wait for Clk_period;
		Addr <=  "0010000010010";
		Trees_din <= x"000b1079";
		wait for Clk_period;
		Addr <=  "0010000010011";
		Trees_din <= x"0203d80c";
		wait for Clk_period;
		Addr <=  "0010000010100";
		Trees_din <= x"08006304";
		wait for Clk_period;
		Addr <=  "0010000010101";
		Trees_din <= x"00381079";
		wait for Clk_period;
		Addr <=  "0010000010110";
		Trees_din <= x"2b009a04";
		wait for Clk_period;
		Addr <=  "0010000010111";
		Trees_din <= x"000b1079";
		wait for Clk_period;
		Addr <=  "0010000011000";
		Trees_din <= x"ff811079";
		wait for Clk_period;
		Addr <=  "0010000011001";
		Trees_din <= x"0d049008";
		wait for Clk_period;
		Addr <=  "0010000011010";
		Trees_din <= x"a807c504";
		wait for Clk_period;
		Addr <=  "0010000011011";
		Trees_din <= x"ffbb1079";
		wait for Clk_period;
		Addr <=  "0010000011100";
		Trees_din <= x"003a1079";
		wait for Clk_period;
		Addr <=  "0010000011101";
		Trees_din <= x"007e1079";
		wait for Clk_period;
		Addr <=  "0010000011110";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0010000011111";
		Trees_din <= x"08016324";
		wait for Clk_period;
		Addr <=  "0010000100000";
		Trees_din <= x"41030b1c";
		wait for Clk_period;
		Addr <=  "0010000100001";
		Trees_din <= x"0d029408";
		wait for Clk_period;
		Addr <=  "0010000100010";
		Trees_din <= x"c608dd04";
		wait for Clk_period;
		Addr <=  "0010000100011";
		Trees_din <= x"ffb11119";
		wait for Clk_period;
		Addr <=  "0010000100100";
		Trees_din <= x"003c1119";
		wait for Clk_period;
		Addr <=  "0010000100101";
		Trees_din <= x"0c03cc0c";
		wait for Clk_period;
		Addr <=  "0010000100110";
		Trees_din <= x"4904ab08";
		wait for Clk_period;
		Addr <=  "0010000100111";
		Trees_din <= x"1605b504";
		wait for Clk_period;
		Addr <=  "0010000101000";
		Trees_din <= x"00961119";
		wait for Clk_period;
		Addr <=  "0010000101001";
		Trees_din <= x"00191119";
		wait for Clk_period;
		Addr <=  "0010000101010";
		Trees_din <= x"fffe1119";
		wait for Clk_period;
		Addr <=  "0010000101011";
		Trees_din <= x"0f04d804";
		wait for Clk_period;
		Addr <=  "0010000101100";
		Trees_din <= x"ffb61119";
		wait for Clk_period;
		Addr <=  "0010000101101";
		Trees_din <= x"003a1119";
		wait for Clk_period;
		Addr <=  "0010000101110";
		Trees_din <= x"2e06f404";
		wait for Clk_period;
		Addr <=  "0010000101111";
		Trees_din <= x"ff961119";
		wait for Clk_period;
		Addr <=  "0010000110000";
		Trees_din <= x"00371119";
		wait for Clk_period;
		Addr <=  "0010000110001";
		Trees_din <= x"0f073b1c";
		wait for Clk_period;
		Addr <=  "0010000110010";
		Trees_din <= x"3501f014";
		wait for Clk_period;
		Addr <=  "0010000110011";
		Trees_din <= x"4f05bc0c";
		wait for Clk_period;
		Addr <=  "0010000110100";
		Trees_din <= x"130a6b08";
		wait for Clk_period;
		Addr <=  "0010000110101";
		Trees_din <= x"ab05eb04";
		wait for Clk_period;
		Addr <=  "0010000110110";
		Trees_din <= x"ff861119";
		wait for Clk_period;
		Addr <=  "0010000110111";
		Trees_din <= x"fff31119";
		wait for Clk_period;
		Addr <=  "0010000111000";
		Trees_din <= x"001a1119";
		wait for Clk_period;
		Addr <=  "0010000111001";
		Trees_din <= x"7400ab04";
		wait for Clk_period;
		Addr <=  "0010000111010";
		Trees_din <= x"00551119";
		wait for Clk_period;
		Addr <=  "0010000111011";
		Trees_din <= x"00141119";
		wait for Clk_period;
		Addr <=  "0010000111100";
		Trees_din <= x"55091b04";
		wait for Clk_period;
		Addr <=  "0010000111101";
		Trees_din <= x"ff6c1119";
		wait for Clk_period;
		Addr <=  "0010000111110";
		Trees_din <= x"fff81119";
		wait for Clk_period;
		Addr <=  "0010000111111";
		Trees_din <= x"1e06630c";
		wait for Clk_period;
		Addr <=  "0010001000000";
		Trees_din <= x"21049108";
		wait for Clk_period;
		Addr <=  "0010001000001";
		Trees_din <= x"03020e04";
		wait for Clk_period;
		Addr <=  "0010001000010";
		Trees_din <= x"fffd1119";
		wait for Clk_period;
		Addr <=  "0010001000011";
		Trees_din <= x"007d1119";
		wait for Clk_period;
		Addr <=  "0010001000100";
		Trees_din <= x"ffd81119";
		wait for Clk_period;
		Addr <=  "0010001000101";
		Trees_din <= x"ffac1119";
		wait for Clk_period;
		Addr <=  "0010001000110";
		Trees_din <= x"12048d2c";
		wait for Clk_period;
		Addr <=  "0010001000111";
		Trees_din <= x"0505e618";
		wait for Clk_period;
		Addr <=  "0010001001000";
		Trees_din <= x"46051208";
		wait for Clk_period;
		Addr <=  "0010001001001";
		Trees_din <= x"dc095e04";
		wait for Clk_period;
		Addr <=  "0010001001010";
		Trees_din <= x"ff6d11ad";
		wait for Clk_period;
		Addr <=  "0010001001011";
		Trees_din <= x"ffcc11ad";
		wait for Clk_period;
		Addr <=  "0010001001100";
		Trees_din <= x"1f03aa04";
		wait for Clk_period;
		Addr <=  "0010001001101";
		Trees_din <= x"ff9511ad";
		wait for Clk_period;
		Addr <=  "0010001001110";
		Trees_din <= x"a9017404";
		wait for Clk_period;
		Addr <=  "0010001001111";
		Trees_din <= x"ffbf11ad";
		wait for Clk_period;
		Addr <=  "0010001010000";
		Trees_din <= x"2303e004";
		wait for Clk_period;
		Addr <=  "0010001010001";
		Trees_din <= x"fffc11ad";
		wait for Clk_period;
		Addr <=  "0010001010010";
		Trees_din <= x"005f11ad";
		wait for Clk_period;
		Addr <=  "0010001010011";
		Trees_din <= x"7401720c";
		wait for Clk_period;
		Addr <=  "0010001010100";
		Trees_din <= x"2e040504";
		wait for Clk_period;
		Addr <=  "0010001010101";
		Trees_din <= x"ffed11ad";
		wait for Clk_period;
		Addr <=  "0010001010110";
		Trees_din <= x"1d021004";
		wait for Clk_period;
		Addr <=  "0010001010111";
		Trees_din <= x"002211ad";
		wait for Clk_period;
		Addr <=  "0010001011000";
		Trees_din <= x"007711ad";
		wait for Clk_period;
		Addr <=  "0010001011001";
		Trees_din <= x"b2008f04";
		wait for Clk_period;
		Addr <=  "0010001011010";
		Trees_din <= x"000511ad";
		wait for Clk_period;
		Addr <=  "0010001011011";
		Trees_din <= x"ff9f11ad";
		wait for Clk_period;
		Addr <=  "0010001011100";
		Trees_din <= x"0904ba18";
		wait for Clk_period;
		Addr <=  "0010001011101";
		Trees_din <= x"16074710";
		wait for Clk_period;
		Addr <=  "0010001011110";
		Trees_din <= x"07050e0c";
		wait for Clk_period;
		Addr <=  "0010001011111";
		Trees_din <= x"0b018404";
		wait for Clk_period;
		Addr <=  "0010001100000";
		Trees_din <= x"ffe511ad";
		wait for Clk_period;
		Addr <=  "0010001100001";
		Trees_din <= x"2b059e04";
		wait for Clk_period;
		Addr <=  "0010001100010";
		Trees_din <= x"008711ad";
		wait for Clk_period;
		Addr <=  "0010001100011";
		Trees_din <= x"000211ad";
		wait for Clk_period;
		Addr <=  "0010001100100";
		Trees_din <= x"ffdb11ad";
		wait for Clk_period;
		Addr <=  "0010001100101";
		Trees_din <= x"1802cc04";
		wait for Clk_period;
		Addr <=  "0010001100110";
		Trees_din <= x"ffab11ad";
		wait for Clk_period;
		Addr <=  "0010001100111";
		Trees_din <= x"fffa11ad";
		wait for Clk_period;
		Addr <=  "0010001101000";
		Trees_din <= x"1502bc04";
		wait for Clk_period;
		Addr <=  "0010001101001";
		Trees_din <= x"001511ad";
		wait for Clk_period;
		Addr <=  "0010001101010";
		Trees_din <= x"ff9411ad";
		wait for Clk_period;
		Addr <=  "0010001101011";
		Trees_din <= x"2c010e28";
		wait for Clk_period;
		Addr <=  "0010001101100";
		Trees_din <= x"56046d18";
		wait for Clk_period;
		Addr <=  "0010001101101";
		Trees_din <= x"ee00db08";
		wait for Clk_period;
		Addr <=  "0010001101110";
		Trees_din <= x"9f05f704";
		wait for Clk_period;
		Addr <=  "0010001101111";
		Trees_din <= x"ffb61239";
		wait for Clk_period;
		Addr <=  "0010001110000";
		Trees_din <= x"003b1239";
		wait for Clk_period;
		Addr <=  "0010001110001";
		Trees_din <= x"8205480c";
		wait for Clk_period;
		Addr <=  "0010001110010";
		Trees_din <= x"4201d704";
		wait for Clk_period;
		Addr <=  "0010001110011";
		Trees_din <= x"fff71239";
		wait for Clk_period;
		Addr <=  "0010001110100";
		Trees_din <= x"3d034304";
		wait for Clk_period;
		Addr <=  "0010001110101";
		Trees_din <= x"008d1239";
		wait for Clk_period;
		Addr <=  "0010001110110";
		Trees_din <= x"00111239";
		wait for Clk_period;
		Addr <=  "0010001110111";
		Trees_din <= x"ffec1239";
		wait for Clk_period;
		Addr <=  "0010001111000";
		Trees_din <= x"03055b0c";
		wait for Clk_period;
		Addr <=  "0010001111001";
		Trees_din <= x"4608fa08";
		wait for Clk_period;
		Addr <=  "0010001111010";
		Trees_din <= x"f0024704";
		wait for Clk_period;
		Addr <=  "0010001111011";
		Trees_din <= x"ff8b1239";
		wait for Clk_period;
		Addr <=  "0010001111100";
		Trees_din <= x"fff61239";
		wait for Clk_period;
		Addr <=  "0010001111101";
		Trees_din <= x"001c1239";
		wait for Clk_period;
		Addr <=  "0010001111110";
		Trees_din <= x"00521239";
		wait for Clk_period;
		Addr <=  "0010001111111";
		Trees_din <= x"1f06af10";
		wait for Clk_period;
		Addr <=  "0010010000000";
		Trees_din <= x"5708b70c";
		wait for Clk_period;
		Addr <=  "0010010000001";
		Trees_din <= x"9c002e04";
		wait for Clk_period;
		Addr <=  "0010010000010";
		Trees_din <= x"fff21239";
		wait for Clk_period;
		Addr <=  "0010010000011";
		Trees_din <= x"19008f04";
		wait for Clk_period;
		Addr <=  "0010010000100";
		Trees_din <= x"ffe01239";
		wait for Clk_period;
		Addr <=  "0010010000101";
		Trees_din <= x"ff701239";
		wait for Clk_period;
		Addr <=  "0010010000110";
		Trees_din <= x"00201239";
		wait for Clk_period;
		Addr <=  "0010010000111";
		Trees_din <= x"0203d808";
		wait for Clk_period;
		Addr <=  "0010010001000";
		Trees_din <= x"2b00fe04";
		wait for Clk_period;
		Addr <=  "0010010001001";
		Trees_din <= x"001b1239";
		wait for Clk_period;
		Addr <=  "0010010001010";
		Trees_din <= x"ffa21239";
		wait for Clk_period;
		Addr <=  "0010010001011";
		Trees_din <= x"66027f04";
		wait for Clk_period;
		Addr <=  "0010010001100";
		Trees_din <= x"fff61239";
		wait for Clk_period;
		Addr <=  "0010010001101";
		Trees_din <= x"00661239";
		wait for Clk_period;
		Addr <=  "0010010001110";
		Trees_din <= x"08013828";
		wait for Clk_period;
		Addr <=  "0010010001111";
		Trees_din <= x"0202dd10";
		wait for Clk_period;
		Addr <=  "0010010010000";
		Trees_din <= x"0b071108";
		wait for Clk_period;
		Addr <=  "0010010010001";
		Trees_din <= x"b800a104";
		wait for Clk_period;
		Addr <=  "0010010010010";
		Trees_din <= x"fff412cd";
		wait for Clk_period;
		Addr <=  "0010010010011";
		Trees_din <= x"ffa112cd";
		wait for Clk_period;
		Addr <=  "0010010010100";
		Trees_din <= x"cc008404";
		wait for Clk_period;
		Addr <=  "0010010010101";
		Trees_din <= x"004312cd";
		wait for Clk_period;
		Addr <=  "0010010010110";
		Trees_din <= x"000312cd";
		wait for Clk_period;
		Addr <=  "0010010010111";
		Trees_din <= x"45026208";
		wait for Clk_period;
		Addr <=  "0010010011000";
		Trees_din <= x"0102d004";
		wait for Clk_period;
		Addr <=  "0010010011001";
		Trees_din <= x"ffb512cd";
		wait for Clk_period;
		Addr <=  "0010010011010";
		Trees_din <= x"003312cd";
		wait for Clk_period;
		Addr <=  "0010010011011";
		Trees_din <= x"3002ef0c";
		wait for Clk_period;
		Addr <=  "0010010011100";
		Trees_din <= x"5606de08";
		wait for Clk_period;
		Addr <=  "0010010011101";
		Trees_din <= x"4c047304";
		wait for Clk_period;
		Addr <=  "0010010011110";
		Trees_din <= x"009112cd";
		wait for Clk_period;
		Addr <=  "0010010011111";
		Trees_din <= x"002712cd";
		wait for Clk_period;
		Addr <=  "0010010100000";
		Trees_din <= x"001012cd";
		wait for Clk_period;
		Addr <=  "0010010100001";
		Trees_din <= x"000c12cd";
		wait for Clk_period;
		Addr <=  "0010010100010";
		Trees_din <= x"0f073b14";
		wait for Clk_period;
		Addr <=  "0010010100011";
		Trees_din <= x"13094a0c";
		wait for Clk_period;
		Addr <=  "0010010100100";
		Trees_din <= x"05097908";
		wait for Clk_period;
		Addr <=  "0010010100101";
		Trees_din <= x"a1096304";
		wait for Clk_period;
		Addr <=  "0010010100110";
		Trees_din <= x"ff7412cd";
		wait for Clk_period;
		Addr <=  "0010010100111";
		Trees_din <= x"ffe212cd";
		wait for Clk_period;
		Addr <=  "0010010101000";
		Trees_din <= x"000712cd";
		wait for Clk_period;
		Addr <=  "0010010101001";
		Trees_din <= x"9f02f604";
		wait for Clk_period;
		Addr <=  "0010010101010";
		Trees_din <= x"ffc412cd";
		wait for Clk_period;
		Addr <=  "0010010101011";
		Trees_din <= x"003e12cd";
		wait for Clk_period;
		Addr <=  "0010010101100";
		Trees_din <= x"4b026a08";
		wait for Clk_period;
		Addr <=  "0010010101101";
		Trees_din <= x"c207d704";
		wait for Clk_period;
		Addr <=  "0010010101110";
		Trees_din <= x"ffad12cd";
		wait for Clk_period;
		Addr <=  "0010010101111";
		Trees_din <= x"000c12cd";
		wait for Clk_period;
		Addr <=  "0010010110000";
		Trees_din <= x"53051804";
		wait for Clk_period;
		Addr <=  "0010010110001";
		Trees_din <= x"007112cd";
		wait for Clk_period;
		Addr <=  "0010010110010";
		Trees_din <= x"fff612cd";
		wait for Clk_period;
		Addr <=  "0010010110011";
		Trees_din <= x"05045024";
		wait for Clk_period;
		Addr <=  "0010010110100";
		Trees_din <= x"8600c918";
		wait for Clk_period;
		Addr <=  "0010010110101";
		Trees_din <= x"08019e0c";
		wait for Clk_period;
		Addr <=  "0010010110110";
		Trees_din <= x"98027c04";
		wait for Clk_period;
		Addr <=  "0010010110111";
		Trees_din <= x"ffe31359";
		wait for Clk_period;
		Addr <=  "0010010111000";
		Trees_din <= x"84020b04";
		wait for Clk_period;
		Addr <=  "0010010111001";
		Trees_din <= x"006e1359";
		wait for Clk_period;
		Addr <=  "0010010111010";
		Trees_din <= x"00181359";
		wait for Clk_period;
		Addr <=  "0010010111011";
		Trees_din <= x"72022108";
		wait for Clk_period;
		Addr <=  "0010010111100";
		Trees_din <= x"95033804";
		wait for Clk_period;
		Addr <=  "0010010111101";
		Trees_din <= x"ffe71359";
		wait for Clk_period;
		Addr <=  "0010010111110";
		Trees_din <= x"ff9e1359";
		wait for Clk_period;
		Addr <=  "0010010111111";
		Trees_din <= x"00191359";
		wait for Clk_period;
		Addr <=  "0010011000000";
		Trees_din <= x"2e076608";
		wait for Clk_period;
		Addr <=  "0010011000001";
		Trees_din <= x"03064904";
		wait for Clk_period;
		Addr <=  "0010011000010";
		Trees_din <= x"ff771359";
		wait for Clk_period;
		Addr <=  "0010011000011";
		Trees_din <= x"ffe21359";
		wait for Clk_period;
		Addr <=  "0010011000100";
		Trees_din <= x"001f1359";
		wait for Clk_period;
		Addr <=  "0010011000101";
		Trees_din <= x"0906421c";
		wait for Clk_period;
		Addr <=  "0010011000110";
		Trees_din <= x"4503ac0c";
		wait for Clk_period;
		Addr <=  "0010011000111";
		Trees_din <= x"0f049004";
		wait for Clk_period;
		Addr <=  "0010011001000";
		Trees_din <= x"ffb01359";
		wait for Clk_period;
		Addr <=  "0010011001001";
		Trees_din <= x"44047604";
		wait for Clk_period;
		Addr <=  "0010011001010";
		Trees_din <= x"fff51359";
		wait for Clk_period;
		Addr <=  "0010011001011";
		Trees_din <= x"00551359";
		wait for Clk_period;
		Addr <=  "0010011001100";
		Trees_din <= x"08035708";
		wait for Clk_period;
		Addr <=  "0010011001101";
		Trees_din <= x"ca002a04";
		wait for Clk_period;
		Addr <=  "0010011001110";
		Trees_din <= x"00131359";
		wait for Clk_period;
		Addr <=  "0010011001111";
		Trees_din <= x"00871359";
		wait for Clk_period;
		Addr <=  "0010011010000";
		Trees_din <= x"ab03de04";
		wait for Clk_period;
		Addr <=  "0010011010001";
		Trees_din <= x"ffe31359";
		wait for Clk_period;
		Addr <=  "0010011010010";
		Trees_din <= x"00441359";
		wait for Clk_period;
		Addr <=  "0010011010011";
		Trees_din <= x"d5015304";
		wait for Clk_period;
		Addr <=  "0010011010100";
		Trees_din <= x"ffa41359";
		wait for Clk_period;
		Addr <=  "0010011010101";
		Trees_din <= x"fff41359";
		wait for Clk_period;
		Addr <=  "0010011010110";
		Trees_din <= x"03041620";
		wait for Clk_period;
		Addr <=  "0010011010111";
		Trees_din <= x"0d04900c";
		wait for Clk_period;
		Addr <=  "0010011011000";
		Trees_din <= x"5507a708";
		wait for Clk_period;
		Addr <=  "0010011011001";
		Trees_din <= x"8200e004";
		wait for Clk_period;
		Addr <=  "0010011011010";
		Trees_din <= x"ffd813cd";
		wait for Clk_period;
		Addr <=  "0010011011011";
		Trees_din <= x"ff7a13cd";
		wait for Clk_period;
		Addr <=  "0010011011100";
		Trees_din <= x"fff513cd";
		wait for Clk_period;
		Addr <=  "0010011011101";
		Trees_din <= x"2303ed08";
		wait for Clk_period;
		Addr <=  "0010011011110";
		Trees_din <= x"c1079904";
		wait for Clk_period;
		Addr <=  "0010011011111";
		Trees_din <= x"ffa613cd";
		wait for Clk_period;
		Addr <=  "0010011100000";
		Trees_din <= x"ffff13cd";
		wait for Clk_period;
		Addr <=  "0010011100001";
		Trees_din <= x"76047108";
		wait for Clk_period;
		Addr <=  "0010011100010";
		Trees_din <= x"0c020b04";
		wait for Clk_period;
		Addr <=  "0010011100011";
		Trees_din <= x"006813cd";
		wait for Clk_period;
		Addr <=  "0010011100100";
		Trees_din <= x"001513cd";
		wait for Clk_period;
		Addr <=  "0010011100101";
		Trees_din <= x"ffdb13cd";
		wait for Clk_period;
		Addr <=  "0010011100110";
		Trees_din <= x"9c01f914";
		wait for Clk_period;
		Addr <=  "0010011100111";
		Trees_din <= x"2f03bf10";
		wait for Clk_period;
		Addr <=  "0010011101000";
		Trees_din <= x"4b025f08";
		wait for Clk_period;
		Addr <=  "0010011101001";
		Trees_din <= x"03080b04";
		wait for Clk_period;
		Addr <=  "0010011101010";
		Trees_din <= x"ffd113cd";
		wait for Clk_period;
		Addr <=  "0010011101011";
		Trees_din <= x"005313cd";
		wait for Clk_period;
		Addr <=  "0010011101100";
		Trees_din <= x"4f023104";
		wait for Clk_period;
		Addr <=  "0010011101101";
		Trees_din <= x"002613cd";
		wait for Clk_period;
		Addr <=  "0010011101110";
		Trees_din <= x"008813cd";
		wait for Clk_period;
		Addr <=  "0010011101111";
		Trees_din <= x"ffe513cd";
		wait for Clk_period;
		Addr <=  "0010011110000";
		Trees_din <= x"39057204";
		wait for Clk_period;
		Addr <=  "0010011110001";
		Trees_din <= x"ffa713cd";
		wait for Clk_period;
		Addr <=  "0010011110010";
		Trees_din <= x"001213cd";
		wait for Clk_period;
		Addr <=  "0010011110011";
		Trees_din <= x"08016c18";
		wait for Clk_period;
		Addr <=  "0010011110100";
		Trees_din <= x"0202dd08";
		wait for Clk_period;
		Addr <=  "0010011110101";
		Trees_din <= x"9c006204";
		wait for Clk_period;
		Addr <=  "0010011110110";
		Trees_din <= x"00271429";
		wait for Clk_period;
		Addr <=  "0010011110111";
		Trees_din <= x"ffb91429";
		wait for Clk_period;
		Addr <=  "0010011111000";
		Trees_din <= x"2301a104";
		wait for Clk_period;
		Addr <=  "0010011111001";
		Trees_din <= x"fff11429";
		wait for Clk_period;
		Addr <=  "0010011111010";
		Trees_din <= x"3002ef08";
		wait for Clk_period;
		Addr <=  "0010011111011";
		Trees_din <= x"76078e04";
		wait for Clk_period;
		Addr <=  "0010011111100";
		Trees_din <= x"00801429";
		wait for Clk_period;
		Addr <=  "0010011111101";
		Trees_din <= x"00151429";
		wait for Clk_period;
		Addr <=  "0010011111110";
		Trees_din <= x"00071429";
		wait for Clk_period;
		Addr <=  "0010011111111";
		Trees_din <= x"5800e010";
		wait for Clk_period;
		Addr <=  "0010100000000";
		Trees_din <= x"4b030208";
		wait for Clk_period;
		Addr <=  "0010100000001";
		Trees_din <= x"18038d04";
		wait for Clk_period;
		Addr <=  "0010100000010";
		Trees_din <= x"ffb41429";
		wait for Clk_period;
		Addr <=  "0010100000011";
		Trees_din <= x"00061429";
		wait for Clk_period;
		Addr <=  "0010100000100";
		Trees_din <= x"6a041a04";
		wait for Clk_period;
		Addr <=  "0010100000101";
		Trees_din <= x"ffea1429";
		wait for Clk_period;
		Addr <=  "0010100000110";
		Trees_din <= x"00551429";
		wait for Clk_period;
		Addr <=  "0010100000111";
		Trees_din <= x"02073404";
		wait for Clk_period;
		Addr <=  "0010100001000";
		Trees_din <= x"ff821429";
		wait for Clk_period;
		Addr <=  "0010100001001";
		Trees_din <= x"fff91429";
		wait for Clk_period;
		Addr <=  "0010100001010";
		Trees_din <= x"0504501c";
		wait for Clk_period;
		Addr <=  "0010100001011";
		Trees_din <= x"8600c910";
		wait for Clk_period;
		Addr <=  "0010100001100";
		Trees_din <= x"0d034204";
		wait for Clk_period;
		Addr <=  "0010100001101";
		Trees_din <= x"ffbe1495";
		wait for Clk_period;
		Addr <=  "0010100001110";
		Trees_din <= x"7505df08";
		wait for Clk_period;
		Addr <=  "0010100001111";
		Trees_din <= x"08019104";
		wait for Clk_period;
		Addr <=  "0010100010000";
		Trees_din <= x"00521495";
		wait for Clk_period;
		Addr <=  "0010100010001";
		Trees_din <= x"00121495";
		wait for Clk_period;
		Addr <=  "0010100010010";
		Trees_din <= x"ffd41495";
		wait for Clk_period;
		Addr <=  "0010100010011";
		Trees_din <= x"2e071308";
		wait for Clk_period;
		Addr <=  "0010100010100";
		Trees_din <= x"1d077804";
		wait for Clk_period;
		Addr <=  "0010100010101";
		Trees_din <= x"ff811495";
		wait for Clk_period;
		Addr <=  "0010100010110";
		Trees_din <= x"ffdd1495";
		wait for Clk_period;
		Addr <=  "0010100010111";
		Trees_din <= x"00151495";
		wait for Clk_period;
		Addr <=  "0010100011000";
		Trees_din <= x"09064218";
		wait for Clk_period;
		Addr <=  "0010100011001";
		Trees_din <= x"4503ac08";
		wait for Clk_period;
		Addr <=  "0010100011010";
		Trees_din <= x"23029f04";
		wait for Clk_period;
		Addr <=  "0010100011011";
		Trees_din <= x"ffc01495";
		wait for Clk_period;
		Addr <=  "0010100011100";
		Trees_din <= x"002a1495";
		wait for Clk_period;
		Addr <=  "0010100011101";
		Trees_din <= x"0301f604";
		wait for Clk_period;
		Addr <=  "0010100011110";
		Trees_din <= x"000f1495";
		wait for Clk_period;
		Addr <=  "0010100011111";
		Trees_din <= x"b8025a08";
		wait for Clk_period;
		Addr <=  "0010100100000";
		Trees_din <= x"8203ed04";
		wait for Clk_period;
		Addr <=  "0010100100001";
		Trees_din <= x"00821495";
		wait for Clk_period;
		Addr <=  "0010100100010";
		Trees_din <= x"00251495";
		wait for Clk_period;
		Addr <=  "0010100100011";
		Trees_din <= x"001c1495";
		wait for Clk_period;
		Addr <=  "0010100100100";
		Trees_din <= x"ffc41495";
		wait for Clk_period;
		Addr <=  "0010100100101";
		Trees_din <= x"2c010e1c";
		wait for Clk_period;
		Addr <=  "0010100100110";
		Trees_din <= x"2e013a0c";
		wait for Clk_period;
		Addr <=  "0010100100111";
		Trees_din <= x"c6070608";
		wait for Clk_period;
		Addr <=  "0010100101000";
		Trees_din <= x"1e043104";
		wait for Clk_period;
		Addr <=  "0010100101001";
		Trees_din <= x"fff314f1";
		wait for Clk_period;
		Addr <=  "0010100101010";
		Trees_din <= x"ffac14f1";
		wait for Clk_period;
		Addr <=  "0010100101011";
		Trees_din <= x"002514f1";
		wait for Clk_period;
		Addr <=  "0010100101100";
		Trees_din <= x"4f01af04";
		wait for Clk_period;
		Addr <=  "0010100101101";
		Trees_din <= x"ffed14f1";
		wait for Clk_period;
		Addr <=  "0010100101110";
		Trees_din <= x"19044b08";
		wait for Clk_period;
		Addr <=  "0010100101111";
		Trees_din <= x"d002aa04";
		wait for Clk_period;
		Addr <=  "0010100110000";
		Trees_din <= x"007c14f1";
		wait for Clk_period;
		Addr <=  "0010100110001";
		Trees_din <= x"002414f1";
		wait for Clk_period;
		Addr <=  "0010100110010";
		Trees_din <= x"fffa14f1";
		wait for Clk_period;
		Addr <=  "0010100110011";
		Trees_din <= x"22013008";
		wait for Clk_period;
		Addr <=  "0010100110100";
		Trees_din <= x"5703cf04";
		wait for Clk_period;
		Addr <=  "0010100110101";
		Trees_din <= x"ffd514f1";
		wait for Clk_period;
		Addr <=  "0010100110110";
		Trees_din <= x"004014f1";
		wait for Clk_period;
		Addr <=  "0010100110111";
		Trees_din <= x"58009808";
		wait for Clk_period;
		Addr <=  "0010100111000";
		Trees_din <= x"8003fa04";
		wait for Clk_period;
		Addr <=  "0010100111001";
		Trees_din <= x"ffd814f1";
		wait for Clk_period;
		Addr <=  "0010100111010";
		Trees_din <= x"001414f1";
		wait for Clk_period;
		Addr <=  "0010100111011";
		Trees_din <= x"ff8614f1";
		wait for Clk_period;
		Addr <=  "0010100111100";
		Trees_din <= x"08013810";
		wait for Clk_period;
		Addr <=  "0010100111101";
		Trees_din <= x"41030b0c";
		wait for Clk_period;
		Addr <=  "0010100111110";
		Trees_din <= x"56045d08";
		wait for Clk_period;
		Addr <=  "0010100111111";
		Trees_din <= x"2c017c04";
		wait for Clk_period;
		Addr <=  "0010101000000";
		Trees_din <= x"0074153d";
		wait for Clk_period;
		Addr <=  "0010101000001";
		Trees_din <= x"0015153d";
		wait for Clk_period;
		Addr <=  "0010101000010";
		Trees_din <= x"fffd153d";
		wait for Clk_period;
		Addr <=  "0010101000011";
		Trees_din <= x"ffdb153d";
		wait for Clk_period;
		Addr <=  "0010101000100";
		Trees_din <= x"6a042908";
		wait for Clk_period;
		Addr <=  "0010101000101";
		Trees_din <= x"4900e304";
		wait for Clk_period;
		Addr <=  "0010101000110";
		Trees_din <= x"ffe7153d";
		wait for Clk_period;
		Addr <=  "0010101000111";
		Trees_din <= x"ff8a153d";
		wait for Clk_period;
		Addr <=  "0010101001000";
		Trees_din <= x"75058608";
		wait for Clk_period;
		Addr <=  "0010101001001";
		Trees_din <= x"f803ed04";
		wait for Clk_period;
		Addr <=  "0010101001010";
		Trees_din <= x"ffe6153d";
		wait for Clk_period;
		Addr <=  "0010101001011";
		Trees_din <= x"004e153d";
		wait for Clk_period;
		Addr <=  "0010101001100";
		Trees_din <= x"f5005204";
		wait for Clk_period;
		Addr <=  "0010101001101";
		Trees_din <= x"fff4153d";
		wait for Clk_period;
		Addr <=  "0010101001110";
		Trees_din <= x"ffaf153d";
		wait for Clk_period;
		Addr <=  "0010101001111";
		Trees_din <= x"03041618";
		wait for Clk_period;
		Addr <=  "0010101010000";
		Trees_din <= x"0d049008";
		wait for Clk_period;
		Addr <=  "0010101010001";
		Trees_din <= x"18049204";
		wait for Clk_period;
		Addr <=  "0010101010010";
		Trees_din <= x"ff911591";
		wait for Clk_period;
		Addr <=  "0010101010011";
		Trees_din <= x"ffe61591";
		wait for Clk_period;
		Addr <=  "0010101010100";
		Trees_din <= x"7a019508";
		wait for Clk_period;
		Addr <=  "0010101010101";
		Trees_din <= x"22015e04";
		wait for Clk_period;
		Addr <=  "0010101010110";
		Trees_din <= x"00431591";
		wait for Clk_period;
		Addr <=  "0010101010111";
		Trees_din <= x"00041591";
		wait for Clk_period;
		Addr <=  "0010101011000";
		Trees_din <= x"92032e04";
		wait for Clk_period;
		Addr <=  "0010101011001";
		Trees_din <= x"fffe1591";
		wait for Clk_period;
		Addr <=  "0010101011010";
		Trees_din <= x"ffbf1591";
		wait for Clk_period;
		Addr <=  "0010101011011";
		Trees_din <= x"1902830c";
		wait for Clk_period;
		Addr <=  "0010101011100";
		Trees_din <= x"0101fb04";
		wait for Clk_period;
		Addr <=  "0010101011101";
		Trees_din <= x"00061591";
		wait for Clk_period;
		Addr <=  "0010101011110";
		Trees_din <= x"75060904";
		wait for Clk_period;
		Addr <=  "0010101011111";
		Trees_din <= x"00751591";
		wait for Clk_period;
		Addr <=  "0010101100000";
		Trees_din <= x"001b1591";
		wait for Clk_period;
		Addr <=  "0010101100001";
		Trees_din <= x"23059404";
		wait for Clk_period;
		Addr <=  "0010101100010";
		Trees_din <= x"ffca1591";
		wait for Clk_period;
		Addr <=  "0010101100011";
		Trees_din <= x"00211591";
		wait for Clk_period;
		Addr <=  "0010101100100";
		Trees_din <= x"05044410";
		wait for Clk_period;
		Addr <=  "0010101100101";
		Trees_din <= x"40009f08";
		wait for Clk_period;
		Addr <=  "0010101100110";
		Trees_din <= x"5602bf04";
		wait for Clk_period;
		Addr <=  "0010101100111";
		Trees_din <= x"003115d5";
		wait for Clk_period;
		Addr <=  "0010101101000";
		Trees_din <= x"ffd515d5";
		wait for Clk_period;
		Addr <=  "0010101101001";
		Trees_din <= x"8600c904";
		wait for Clk_period;
		Addr <=  "0010101101010";
		Trees_din <= x"ffee15d5";
		wait for Clk_period;
		Addr <=  "0010101101011";
		Trees_din <= x"ff9715d5";
		wait for Clk_period;
		Addr <=  "0010101101100";
		Trees_din <= x"b1018e04";
		wait for Clk_period;
		Addr <=  "0010101101101";
		Trees_din <= x"ffd015d5";
		wait for Clk_period;
		Addr <=  "0010101101110";
		Trees_din <= x"2b04e40c";
		wait for Clk_period;
		Addr <=  "0010101101111";
		Trees_din <= x"07045608";
		wait for Clk_period;
		Addr <=  "0010101110000";
		Trees_din <= x"21042004";
		wait for Clk_period;
		Addr <=  "0010101110001";
		Trees_din <= x"007015d5";
		wait for Clk_period;
		Addr <=  "0010101110010";
		Trees_din <= x"001715d5";
		wait for Clk_period;
		Addr <=  "0010101110011";
		Trees_din <= x"fffa15d5";
		wait for Clk_period;
		Addr <=  "0010101110100";
		Trees_din <= x"ffec15d5";
		wait for Clk_period;
		Addr <=  "0010101110101";
		Trees_din <= x"08019e10";
		wait for Clk_period;
		Addr <=  "0010101110110";
		Trees_din <= x"02026404";
		wait for Clk_period;
		Addr <=  "0010101110111";
		Trees_din <= x"ffde1619";
		wait for Clk_period;
		Addr <=  "0010101111000";
		Trees_din <= x"b3026708";
		wait for Clk_period;
		Addr <=  "0010101111001";
		Trees_din <= x"43032e04";
		wait for Clk_period;
		Addr <=  "0010101111010";
		Trees_din <= x"00661619";
		wait for Clk_period;
		Addr <=  "0010101111011";
		Trees_din <= x"00171619";
		wait for Clk_period;
		Addr <=  "0010101111100";
		Trees_din <= x"fff21619";
		wait for Clk_period;
		Addr <=  "0010101111101";
		Trees_din <= x"5800980c";
		wait for Clk_period;
		Addr <=  "0010101111110";
		Trees_din <= x"1e04af08";
		wait for Clk_period;
		Addr <=  "0010101111111";
		Trees_din <= x"4e05a304";
		wait for Clk_period;
		Addr <=  "0010110000000";
		Trees_din <= x"fff21619";
		wait for Clk_period;
		Addr <=  "0010110000001";
		Trees_din <= x"00431619";
		wait for Clk_period;
		Addr <=  "0010110000010";
		Trees_din <= x"ffd11619";
		wait for Clk_period;
		Addr <=  "0010110000011";
		Trees_din <= x"bd059304";
		wait for Clk_period;
		Addr <=  "0010110000100";
		Trees_din <= x"ff961619";
		wait for Clk_period;
		Addr <=  "0010110000101";
		Trees_din <= x"ffef1619";
		wait for Clk_period;
		Addr <=  "0010110000110";
		Trees_din <= x"02056014";
		wait for Clk_period;
		Addr <=  "0010110000111";
		Trees_din <= x"0d04a108";
		wait for Clk_period;
		Addr <=  "0010110001000";
		Trees_din <= x"0b06e604";
		wait for Clk_period;
		Addr <=  "0010110001001";
		Trees_din <= x"ff9b1655";
		wait for Clk_period;
		Addr <=  "0010110001010";
		Trees_din <= x"fff91655";
		wait for Clk_period;
		Addr <=  "0010110001011";
		Trees_din <= x"22027208";
		wait for Clk_period;
		Addr <=  "0010110001100";
		Trees_din <= x"4203bc04";
		wait for Clk_period;
		Addr <=  "0010110001101";
		Trees_din <= x"fff91655";
		wait for Clk_period;
		Addr <=  "0010110001110";
		Trees_din <= x"00431655";
		wait for Clk_period;
		Addr <=  "0010110001111";
		Trees_din <= x"ffcd1655";
		wait for Clk_period;
		Addr <=  "0010110010000";
		Trees_din <= x"2104e708";
		wait for Clk_period;
		Addr <=  "0010110010001";
		Trees_din <= x"07029604";
		wait for Clk_period;
		Addr <=  "0010110010010";
		Trees_din <= x"00611655";
		wait for Clk_period;
		Addr <=  "0010110010011";
		Trees_din <= x"00071655";
		wait for Clk_period;
		Addr <=  "0010110010100";
		Trees_din <= x"ffeb1655";
		wait for Clk_period;
		Addr <=  "0010110010101";
		Trees_din <= x"1203510c";
		wait for Clk_period;
		Addr <=  "0010110010110";
		Trees_din <= x"0506b608";
		wait for Clk_period;
		Addr <=  "0010110010111";
		Trees_din <= x"3a00f904";
		wait for Clk_period;
		Addr <=  "0010110011000";
		Trees_din <= x"ffe91691";
		wait for Clk_period;
		Addr <=  "0010110011001";
		Trees_din <= x"ff9f1691";
		wait for Clk_period;
		Addr <=  "0010110011010";
		Trees_din <= x"00051691";
		wait for Clk_period;
		Addr <=  "0010110011011";
		Trees_din <= x"0304160c";
		wait for Clk_period;
		Addr <=  "0010110011100";
		Trees_din <= x"a104fd08";
		wait for Clk_period;
		Addr <=  "0010110011101";
		Trees_din <= x"0a02b204";
		wait for Clk_period;
		Addr <=  "0010110011110";
		Trees_din <= x"fff81691";
		wait for Clk_period;
		Addr <=  "0010110011111";
		Trees_din <= x"ffbf1691";
		wait for Clk_period;
		Addr <=  "0010110100000";
		Trees_din <= x"00221691";
		wait for Clk_period;
		Addr <=  "0010110100001";
		Trees_din <= x"39035d04";
		wait for Clk_period;
		Addr <=  "0010110100010";
		Trees_din <= x"fff71691";
		wait for Clk_period;
		Addr <=  "0010110100011";
		Trees_din <= x"005d1691";
		wait for Clk_period;
		Addr <=  "0010110100100";
		Trees_din <= x"0f069314";
		wait for Clk_period;
		Addr <=  "0010110100101";
		Trees_din <= x"c701070c";
		wait for Clk_period;
		Addr <=  "0010110100110";
		Trees_din <= x"5301ff08";
		wait for Clk_period;
		Addr <=  "0010110100111";
		Trees_din <= x"2e042a04";
		wait for Clk_period;
		Addr <=  "0010110101000";
		Trees_din <= x"000f16cd";
		wait for Clk_period;
		Addr <=  "0010110101001";
		Trees_din <= x"003a16cd";
		wait for Clk_period;
		Addr <=  "0010110101010";
		Trees_din <= x"ffdc16cd";
		wait for Clk_period;
		Addr <=  "0010110101011";
		Trees_din <= x"7800e204";
		wait for Clk_period;
		Addr <=  "0010110101100";
		Trees_din <= x"fff816cd";
		wait for Clk_period;
		Addr <=  "0010110101101";
		Trees_din <= x"ffa816cd";
		wait for Clk_period;
		Addr <=  "0010110101110";
		Trees_din <= x"2e00d804";
		wait for Clk_period;
		Addr <=  "0010110101111";
		Trees_din <= x"fff116cd";
		wait for Clk_period;
		Addr <=  "0010110110000";
		Trees_din <= x"4603a304";
		wait for Clk_period;
		Addr <=  "0010110110001";
		Trees_din <= x"001916cd";
		wait for Clk_period;
		Addr <=  "0010110110010";
		Trees_din <= x"005d16cd";
		wait for Clk_period;
		Addr <=  "0010110110011";
		Trees_din <= x"08016c0c";
		wait for Clk_period;
		Addr <=  "0010110110100";
		Trees_din <= x"14033e08";
		wait for Clk_period;
		Addr <=  "0010110110101";
		Trees_din <= x"7b025704";
		wait for Clk_period;
		Addr <=  "0010110110110";
		Trees_din <= x"00541701";
		wait for Clk_period;
		Addr <=  "0010110110111";
		Trees_din <= x"00011701";
		wait for Clk_period;
		Addr <=  "0010110111000";
		Trees_din <= x"fff01701";
		wait for Clk_period;
		Addr <=  "0010110111001";
		Trees_din <= x"58009808";
		wait for Clk_period;
		Addr <=  "0010110111010";
		Trees_din <= x"4b032b04";
		wait for Clk_period;
		Addr <=  "0010110111011";
		Trees_din <= x"ffe51701";
		wait for Clk_period;
		Addr <=  "0010110111100";
		Trees_din <= x"00271701";
		wait for Clk_period;
		Addr <=  "0010110111101";
		Trees_din <= x"0105c604";
		wait for Clk_period;
		Addr <=  "0010110111110";
		Trees_din <= x"ffa81701";
		wait for Clk_period;
		Addr <=  "0010110111111";
		Trees_din <= x"ffec1701";
		wait for Clk_period;
		Addr <=  "0010111000000";
		Trees_din <= x"0503c50c";
		wait for Clk_period;
		Addr <=  "0010111000001";
		Trees_din <= x"9b058408";
		wait for Clk_period;
		Addr <=  "0010111000010";
		Trees_din <= x"34052804";
		wait for Clk_period;
		Addr <=  "0010111000011";
		Trees_din <= x"ffac1735";
		wait for Clk_period;
		Addr <=  "0010111000100";
		Trees_din <= x"fff01735";
		wait for Clk_period;
		Addr <=  "0010111000101";
		Trees_din <= x"00091735";
		wait for Clk_period;
		Addr <=  "0010111000110";
		Trees_din <= x"1903490c";
		wait for Clk_period;
		Addr <=  "0010111000111";
		Trees_din <= x"12037b04";
		wait for Clk_period;
		Addr <=  "0010111001000";
		Trees_din <= x"fffe1735";
		wait for Clk_period;
		Addr <=  "0010111001001";
		Trees_din <= x"18022f04";
		wait for Clk_period;
		Addr <=  "0010111001010";
		Trees_din <= x"00101735";
		wait for Clk_period;
		Addr <=  "0010111001011";
		Trees_din <= x"005d1735";
		wait for Clk_period;
		Addr <=  "0010111001100";
		Trees_din <= x"ffe61735";
		wait for Clk_period;
		Addr <=  "0010111001101";
		Trees_din <= x"e4022810";
		wait for Clk_period;
		Addr <=  "0010111001110";
		Trees_din <= x"2301a104";
		wait for Clk_period;
		Addr <=  "0010111001111";
		Trees_din <= x"ffd31761";
		wait for Clk_period;
		Addr <=  "0010111010000";
		Trees_din <= x"8203ed08";
		wait for Clk_period;
		Addr <=  "0010111010001";
		Trees_din <= x"8a028304";
		wait for Clk_period;
		Addr <=  "0010111010010";
		Trees_din <= x"00591761";
		wait for Clk_period;
		Addr <=  "0010111010011";
		Trees_din <= x"000b1761";
		wait for Clk_period;
		Addr <=  "0010111010100";
		Trees_din <= x"ffe91761";
		wait for Clk_period;
		Addr <=  "0010111010101";
		Trees_din <= x"18046404";
		wait for Clk_period;
		Addr <=  "0010111010110";
		Trees_din <= x"ffb01761";
		wait for Clk_period;
		Addr <=  "0010111010111";
		Trees_din <= x"00041761";
		wait for Clk_period;
		Addr <=  "0010111011000";
		Trees_din <= x"2c00e810";
		wait for Clk_period;
		Addr <=  "0010111011001";
		Trees_din <= x"7904e60c";
		wait for Clk_period;
		Addr <=  "0010111011010";
		Trees_din <= x"16035708";
		wait for Clk_period;
		Addr <=  "0010111011011";
		Trees_din <= x"39044704";
		wait for Clk_period;
		Addr <=  "0010111011100";
		Trees_din <= x"00101795";
		wait for Clk_period;
		Addr <=  "0010111011101";
		Trees_din <= x"00581795";
		wait for Clk_period;
		Addr <=  "0010111011110";
		Trees_din <= x"fffc1795";
		wait for Clk_period;
		Addr <=  "0010111011111";
		Trees_din <= x"ffdd1795";
		wait for Clk_period;
		Addr <=  "0010111100000";
		Trees_din <= x"13079008";
		wait for Clk_period;
		Addr <=  "0010111100001";
		Trees_din <= x"2303ed04";
		wait for Clk_period;
		Addr <=  "0010111100010";
		Trees_din <= x"ffab1795";
		wait for Clk_period;
		Addr <=  "0010111100011";
		Trees_din <= x"ffeb1795";
		wait for Clk_period;
		Addr <=  "0010111100100";
		Trees_din <= x"00141795";
		wait for Clk_period;
		Addr <=  "0010111100101";
		Trees_din <= x"2e04320c";
		wait for Clk_period;
		Addr <=  "0010111100110";
		Trees_din <= x"1206ef08";
		wait for Clk_period;
		Addr <=  "0010111100111";
		Trees_din <= x"1804ed04";
		wait for Clk_period;
		Addr <=  "0010111101000";
		Trees_din <= x"ffb117b9";
		wait for Clk_period;
		Addr <=  "0010111101001";
		Trees_din <= x"fffc17b9";
		wait for Clk_period;
		Addr <=  "0010111101010";
		Trees_din <= x"001517b9";
		wait for Clk_period;
		Addr <=  "0010111101011";
		Trees_din <= x"0f031d04";
		wait for Clk_period;
		Addr <=  "0010111101100";
		Trees_din <= x"fff417b9";
		wait for Clk_period;
		Addr <=  "0010111101101";
		Trees_din <= x"004417b9";
		wait for Clk_period;
		Addr <=  "0010111101110";
		Trees_din <= x"0801380c";
		wait for Clk_period;
		Addr <=  "0010111101111";
		Trees_din <= x"2c016908";
		wait for Clk_period;
		Addr <=  "0010111110000";
		Trees_din <= x"9802fe04";
		wait for Clk_period;
		Addr <=  "0010111110001";
		Trees_din <= x"000617e5";
		wait for Clk_period;
		Addr <=  "0010111110010";
		Trees_din <= x"004817e5";
		wait for Clk_period;
		Addr <=  "0010111110011";
		Trees_din <= x"fff017e5";
		wait for Clk_period;
		Addr <=  "0010111110100";
		Trees_din <= x"2100ce04";
		wait for Clk_period;
		Addr <=  "0010111110101";
		Trees_din <= x"001317e5";
		wait for Clk_period;
		Addr <=  "0010111110110";
		Trees_din <= x"18052b04";
		wait for Clk_period;
		Addr <=  "0010111110111";
		Trees_din <= x"ffb217e5";
		wait for Clk_period;
		Addr <=  "0010111111000";
		Trees_din <= x"fffe17e5";
		wait for Clk_period;
		Addr <=  "0010111111001";
		Trees_din <= x"0205600c";
		wait for Clk_period;
		Addr <=  "0010111111010";
		Trees_din <= x"83007204";
		wait for Clk_period;
		Addr <=  "0010111111011";
		Trees_din <= x"000f1809";
		wait for Clk_period;
		Addr <=  "0010111111100";
		Trees_din <= x"5d05c804";
		wait for Clk_period;
		Addr <=  "0010111111101";
		Trees_din <= x"ffb51809";
		wait for Clk_period;
		Addr <=  "0010111111110";
		Trees_din <= x"fff21809";
		wait for Clk_period;
		Addr <=  "0010111111111";
		Trees_din <= x"2e03fc04";
		wait for Clk_period;
		Addr <=  "0011000000000";
		Trees_din <= x"fffe1809";
		wait for Clk_period;
		Addr <=  "0011000000001";
		Trees_din <= x"00421809";
		wait for Clk_period;
		Addr <=  "0011000000010";
		Trees_din <= x"05073b10";
		wait for Clk_period;
		Addr <=  "0011000000011";
		Trees_din <= x"53020308";
		wait for Clk_period;
		Addr <=  "0011000000100";
		Trees_din <= x"1d03e304";
		wait for Clk_period;
		Addr <=  "0011000000101";
		Trees_din <= x"ffe91835";
		wait for Clk_period;
		Addr <=  "0011000000110";
		Trees_din <= x"00271835";
		wait for Clk_period;
		Addr <=  "0011000000111";
		Trees_din <= x"0d063904";
		wait for Clk_period;
		Addr <=  "0011000001000";
		Trees_din <= x"ffb81835";
		wait for Clk_period;
		Addr <=  "0011000001001";
		Trees_din <= x"fffd1835";
		wait for Clk_period;
		Addr <=  "0011000001010";
		Trees_din <= x"1803a804";
		wait for Clk_period;
		Addr <=  "0011000001011";
		Trees_din <= x"00071835";
		wait for Clk_period;
		Addr <=  "0011000001100";
		Trees_din <= x"00411835";
		wait for Clk_period;
		Addr <=  "0011000001101";
		Trees_din <= x"02026408";
		wait for Clk_period;
		Addr <=  "0011000001110";
		Trees_din <= x"34053704";
		wait for Clk_period;
		Addr <=  "0011000001111";
		Trees_din <= x"ffbd1859";
		wait for Clk_period;
		Addr <=  "0011000010000";
		Trees_din <= x"fffd1859";
		wait for Clk_period;
		Addr <=  "0011000010001";
		Trees_din <= x"21040d08";
		wait for Clk_period;
		Addr <=  "0011000010010";
		Trees_din <= x"0801c504";
		wait for Clk_period;
		Addr <=  "0011000010011";
		Trees_din <= x"003f1859";
		wait for Clk_period;
		Addr <=  "0011000010100";
		Trees_din <= x"fffe1859";
		wait for Clk_period;
		Addr <=  "0011000010101";
		Trees_din <= x"ffe41859";
		wait for Clk_period;
		Addr <=  "0011000010110";
		Trees_din <= x"0f06930c";
		wait for Clk_period;
		Addr <=  "0011000010111";
		Trees_din <= x"f1011308";
		wait for Clk_period;
		Addr <=  "0011000011000";
		Trees_din <= x"b8016704";
		wait for Clk_period;
		Addr <=  "0011000011001";
		Trees_din <= x"0028187d";
		wait for Clk_period;
		Addr <=  "0011000011010";
		Trees_din <= x"ffeb187d";
		wait for Clk_period;
		Addr <=  "0011000011011";
		Trees_din <= x"ffc3187d";
		wait for Clk_period;
		Addr <=  "0011000011100";
		Trees_din <= x"4604d204";
		wait for Clk_period;
		Addr <=  "0011000011101";
		Trees_din <= x"fffa187d";
		wait for Clk_period;
		Addr <=  "0011000011110";
		Trees_din <= x"0042187d";
		wait for Clk_period;
		Addr <=  "0011000011111";
		Trees_din <= x"2c00e80c";
		wait for Clk_period;
		Addr <=  "0011000100000";
		Trees_din <= x"4b020e04";
		wait for Clk_period;
		Addr <=  "0011000100001";
		Trees_din <= x"ffed18a1";
		wait for Clk_period;
		Addr <=  "0011000100010";
		Trees_din <= x"9f03c004";
		wait for Clk_period;
		Addr <=  "0011000100011";
		Trees_din <= x"000e18a1";
		wait for Clk_period;
		Addr <=  "0011000100100";
		Trees_din <= x"004318a1";
		wait for Clk_period;
		Addr <=  "0011000100101";
		Trees_din <= x"0203d804";
		wait for Clk_period;
		Addr <=  "0011000100110";
		Trees_din <= x"ffc518a1";
		wait for Clk_period;
		Addr <=  "0011000100111";
		Trees_din <= x"000118a1";
		wait for Clk_period;
		Addr <=  "0011000101000";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  5
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"360b8c30";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"11112c24";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"2112a11c";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"0100000c";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"4c01fd08";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"4b023504";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"02240095";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"ff750095";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"ff560095";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"3607b408";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"110cfd04";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"ff4e0095";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"ff890095";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"7906e704";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"ff5e0095";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"00400095";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"01012e04";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"013c0095";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"ff850095";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"2109e008";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"1605fb04";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"ff620095";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"00b20095";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"02e40095";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"2104a60c";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"38007904";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"01640095";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"13015b04";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"00270095";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"ff590095";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"34052808";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"27032204";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"00270095";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"038b0095";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"0201e204";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"00b20095";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"ff810095";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"360afc30";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"2112a128";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"11134620";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"2706df10";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"97000108";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"70008104";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"ff770139";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"00ca0139";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"400d4d04";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"ff550139";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"ffef0139";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"ca066308";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"3605cc04";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"ff9a0139";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"01710139";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"6405c804";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"ff5a0139";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"001f0139";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"05054504";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"01660139";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"ff840139";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"79094e04";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"ff880139";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"01980139";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"45051318";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"0c045d10";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"6c07be0c";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"7d028608";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"31086f04";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"020f0139";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"00930139";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"ff9d0139";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"ff970139";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"14020204";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"00bb0139";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"ff740139";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"1c094b04";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"ff5d0139";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"1f00a904";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"011e0139";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"00320139";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"360afc30";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"2112a128";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"11134620";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"2706df10";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"97000108";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"0a023c04";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"00d401d5";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"ff7d01d5";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"1b0ee404";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"ff5a01d5";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"000101d5";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"6c00c008";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"0202a704";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"ff8701d5";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"01a401d5";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"5804b504";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"ff5f01d5";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"000701d5";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"05054504";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"011401d5";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"ff8e01d5";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"1b063104";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"ff9001d5";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"013001d5";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"0d049018";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"f901f510";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"83007604";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"ff9901d5";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"3c080c08";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"5000d204";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"000301d5";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"015701d5";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"ffa601d5";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"35094404";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"ff7c01d5";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"002501d5";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"4a033e04";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"ff6601d5";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"002601d5";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"360afc3c";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"110ec730";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"3607b41c";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"0100000c";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"2105f004";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"ff6a0291";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"ab018d04";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"013c0291";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"ff9f0291";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"720b6a08";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"110cfd04";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"ff5e0291";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"ffb90291";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"d602f704";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"00450291";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"ffa90291";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"7906e708";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"b3051204";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"ff600291";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"005e0291";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"d7031908";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"d2040104";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"ffa80291";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"016a0291";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"ff840291";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"4006e604";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"ff6a0291";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"0d033a04";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"01550291";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"fff70291";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"4505131c";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"1b02a308";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"bc030b04";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"00110291";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"ff8a0291";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"bb002004";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"ffa20291";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"13080808";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"ce07f304";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"01240291";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"00580291";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"1500a604";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"ffaa0291";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"006d0291";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"1c094b04";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"ff680291";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"00a00291";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"360afc2c";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"110ec720";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"ba073510";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"3e14d20c";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"11085f04";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"ff5f0325";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"45008404";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"00830325";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"ff6d0325";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"00160325";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"3001d204";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"ff600325";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"11047b04";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"ff6b0325";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"01036504";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"013e0325";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"ff810325";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"4006e604";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"ff700325";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"0d033a04";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"01130325";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"fffa0325";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"0d049018";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"4d040308";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"1b04ee04";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"ff800325";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"007d0325";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"6800a604";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"ffaa0325";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"48034c08";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"7d019c04";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"00f60325";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"00540325";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"00200325";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"e50d0504";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"ff730325";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"000c0325";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"3608b238";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"110cfd24";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"0100000c";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"2105f004";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"ff7603d1";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"4c01fd04";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"00cf03d1";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"ffad03d1";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"a50c7d10";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"1c0a1a08";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"520c8e04";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"ff6303d1";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"000a03d1";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"1700b504";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"009303d1";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"ff8703d1";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"4e00b004";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"00b903d1";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"ff9203d1";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"0d03f70c";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"83039004";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"ff9f03d1";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"5b005504";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"003b03d1";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"011b03d1";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"12011f04";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"001803d1";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"ff7003d1";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"0d03f718";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"11042e04";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"ff8403d1";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"09016c0c";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"6b030504";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"ffa703d1";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"1c00ef04";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"ffd803d1";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"00de03d1";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"de004004";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"004603d1";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"ff8b03d1";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"38005504";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"004503d1";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"ff6a03d1";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"3608b240";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"11068820";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"b20b5318";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"05000608";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"3d013004";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"00440495";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"ff8c0495";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"b7000108";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"b2050f04";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"ff7f0495";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"004a0495";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"08000004";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"ffb80495";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"ff620495";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"4d004604";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"00320495";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"ffb00495";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"0101c710";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"ae02520c";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"5b039008";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"8d00b504";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"ffe00495";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"01230495";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"ff890495";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"ff760495";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"8605d608";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"11134604";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"ff650495";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"00080495";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"dc068504";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"ffaa0495";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"00910495";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"0d041e1c";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"11042e04";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"ff8a0495";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"09016c10";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"4505d308";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"4d025004";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"ffef0495";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"00cf0495";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"97000704";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"00800495";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"ff930495";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"7f009304";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"00380495";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"ff940495";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"350bc404";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"ff6e0495";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"003c0495";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"1b074b44";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"27067118";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"97000108";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"0e00e104";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"00790565";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"ffac0565";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"400c530c";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"b7000108";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"5f019504";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"ff8c0565";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"004a0565";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"ff630565";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"00240565";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"d7031d18";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"4a00db0c";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"f8015a04";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"008e0565";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"13018e04";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"fff40565";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"ff7d0565";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"1f052508";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"0101c704";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"00fd0565";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"002b0565";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"00010565";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"6c02be0c";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"d0057908";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"98014d04";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"ffea0565";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"ff8e0565";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"007a0565";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"46007c04";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"ffd80565";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"ff680565";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"0d025d14";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"6b030e04";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"ff940565";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"1d05a50c";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"01068d08";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"29045804";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"00da0565";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"003f0565";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"001a0565";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"ffbf0565";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"aa048d0c";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"210cb808";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"70000004";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"fff00565";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"ff6e0565";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"00240565";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"00950565";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"1b074b34";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"27067114";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"97000104";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"00160611";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"400c530c";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"b7000108";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"dd061d04";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"ff950611";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"004b0611";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"ff640611";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"00210611";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"d7031d10";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"3405720c";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"1f05cb08";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"80026c04";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"00040611";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"00dd0611";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"ffa40611";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"ff8a0611";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"d0067c08";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"3b096204";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"ff6a0611";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"00050611";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"96025304";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"ff9c0611";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"007b0611";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"0d025d14";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"6b030e04";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"ff9d0611";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"1d05a50c";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"58000504";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"00110611";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"3a01df04";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"00cc0611";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"003f0611";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"ffc70611";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"aa048d0c";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"210cb808";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"26000404";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"ffed0611";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"ff720611";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"00200611";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"00850611";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"1b074b34";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"27067114";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"97000104";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"001506b5";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"400c530c";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"b7000108";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"f3058204";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"ff9e06b5";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"004b06b5";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"ff6506b5";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"001c06b5";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"d7031d10";
		wait for Clk_period;
		Addr <=  "0000110010000";
		Trees_din <= x"3405720c";
		wait for Clk_period;
		Addr <=  "0000110010001";
		Trees_din <= x"1f05cb08";
		wait for Clk_period;
		Addr <=  "0000110010010";
		Trees_din <= x"80026c04";
		wait for Clk_period;
		Addr <=  "0000110010011";
		Trees_din <= x"000406b5";
		wait for Clk_period;
		Addr <=  "0000110010100";
		Trees_din <= x"00c406b5";
		wait for Clk_period;
		Addr <=  "0000110010101";
		Trees_din <= x"ffac06b5";
		wait for Clk_period;
		Addr <=  "0000110010110";
		Trees_din <= x"ff9206b5";
		wait for Clk_period;
		Addr <=  "0000110010111";
		Trees_din <= x"92059d08";
		wait for Clk_period;
		Addr <=  "0000110011000";
		Trees_din <= x"4a032004";
		wait for Clk_period;
		Addr <=  "0000110011001";
		Trees_din <= x"ff6d06b5";
		wait for Clk_period;
		Addr <=  "0000110011010";
		Trees_din <= x"ffea06b5";
		wait for Clk_period;
		Addr <=  "0000110011011";
		Trees_din <= x"6c02be04";
		wait for Clk_period;
		Addr <=  "0000110011100";
		Trees_din <= x"005e06b5";
		wait for Clk_period;
		Addr <=  "0000110011101";
		Trees_din <= x"ffb806b5";
		wait for Clk_period;
		Addr <=  "0000110011110";
		Trees_din <= x"c2018e0c";
		wait for Clk_period;
		Addr <=  "0000110011111";
		Trees_din <= x"4d03ec04";
		wait for Clk_period;
		Addr <=  "0000110100000";
		Trees_din <= x"ffb106b5";
		wait for Clk_period;
		Addr <=  "0000110100001";
		Trees_din <= x"f900cc04";
		wait for Clk_period;
		Addr <=  "0000110100010";
		Trees_din <= x"00c806b5";
		wait for Clk_period;
		Addr <=  "0000110100011";
		Trees_din <= x"001b06b5";
		wait for Clk_period;
		Addr <=  "0000110100100";
		Trees_din <= x"21051004";
		wait for Clk_period;
		Addr <=  "0000110100101";
		Trees_din <= x"ff7d06b5";
		wait for Clk_period;
		Addr <=  "0000110100110";
		Trees_din <= x"2705d808";
		wait for Clk_period;
		Addr <=  "0000110100111";
		Trees_din <= x"c5003804";
		wait for Clk_period;
		Addr <=  "0000110101000";
		Trees_din <= x"000806b5";
		wait for Clk_period;
		Addr <=  "0000110101001";
		Trees_din <= x"ff9c06b5";
		wait for Clk_period;
		Addr <=  "0000110101010";
		Trees_din <= x"80013904";
		wait for Clk_period;
		Addr <=  "0000110101011";
		Trees_din <= x"002306b5";
		wait for Clk_period;
		Addr <=  "0000110101100";
		Trees_din <= x"009606b5";
		wait for Clk_period;
		Addr <=  "0000110101101";
		Trees_din <= x"ba073524";
		wait for Clk_period;
		Addr <=  "0000110101110";
		Trees_din <= x"400c531c";
		wait for Clk_period;
		Addr <=  "0000110101111";
		Trees_din <= x"11082d10";
		wait for Clk_period;
		Addr <=  "0000110110000";
		Trees_din <= x"b7000108";
		wait for Clk_period;
		Addr <=  "0000110110001";
		Trees_din <= x"1201c804";
		wait for Clk_period;
		Addr <=  "0000110110010";
		Trees_din <= x"004b0739";
		wait for Clk_period;
		Addr <=  "0000110110011";
		Trees_din <= x"ffa30739";
		wait for Clk_period;
		Addr <=  "0000110110100";
		Trees_din <= x"720a4704";
		wait for Clk_period;
		Addr <=  "0000110110101";
		Trees_din <= x"ff660739";
		wait for Clk_period;
		Addr <=  "0000110110110";
		Trees_din <= x"ffee0739";
		wait for Clk_period;
		Addr <=  "0000110110111";
		Trees_din <= x"c8002504";
		wait for Clk_period;
		Addr <=  "0000110111000";
		Trees_din <= x"00820739";
		wait for Clk_period;
		Addr <=  "0000110111001";
		Trees_din <= x"30052404";
		wait for Clk_period;
		Addr <=  "0000110111010";
		Trees_din <= x"ff750739";
		wait for Clk_period;
		Addr <=  "0000110111011";
		Trees_din <= x"00240739";
		wait for Clk_period;
		Addr <=  "0000110111100";
		Trees_din <= x"97035904";
		wait for Clk_period;
		Addr <=  "0000110111101";
		Trees_din <= x"ffd90739";
		wait for Clk_period;
		Addr <=  "0000110111110";
		Trees_din <= x"00620739";
		wait for Clk_period;
		Addr <=  "0000110111111";
		Trees_din <= x"3404b818";
		wait for Clk_period;
		Addr <=  "0000111000000";
		Trees_din <= x"6400c208";
		wait for Clk_period;
		Addr <=  "0000111000001";
		Trees_din <= x"1c06a304";
		wait for Clk_period;
		Addr <=  "0000111000010";
		Trees_din <= x"ff850739";
		wait for Clk_period;
		Addr <=  "0000111000011";
		Trees_din <= x"002c0739";
		wait for Clk_period;
		Addr <=  "0000111000100";
		Trees_din <= x"11042e04";
		wait for Clk_period;
		Addr <=  "0000111000101";
		Trees_din <= x"ffb10739";
		wait for Clk_period;
		Addr <=  "0000111000110";
		Trees_din <= x"41036a08";
		wait for Clk_period;
		Addr <=  "0000111000111";
		Trees_din <= x"1c021d04";
		wait for Clk_period;
		Addr <=  "0000111001000";
		Trees_din <= x"001c0739";
		wait for Clk_period;
		Addr <=  "0000111001001";
		Trees_din <= x"00b40739";
		wait for Clk_period;
		Addr <=  "0000111001010";
		Trees_din <= x"ffd70739";
		wait for Clk_period;
		Addr <=  "0000111001011";
		Trees_din <= x"17000004";
		wait for Clk_period;
		Addr <=  "0000111001100";
		Trees_din <= x"fffc0739";
		wait for Clk_period;
		Addr <=  "0000111001101";
		Trees_din <= x"ff700739";
		wait for Clk_period;
		Addr <=  "0000111001110";
		Trees_din <= x"1b074b30";
		wait for Clk_period;
		Addr <=  "0000111001111";
		Trees_din <= x"27067114";
		wait for Clk_period;
		Addr <=  "0000111010000";
		Trees_din <= x"97000104";
		wait for Clk_period;
		Addr <=  "0000111010001";
		Trees_din <= x"001907cd";
		wait for Clk_period;
		Addr <=  "0000111010010";
		Trees_din <= x"b7000108";
		wait for Clk_period;
		Addr <=  "0000111010011";
		Trees_din <= x"49021c04";
		wait for Clk_period;
		Addr <=  "0000111010100";
		Trees_din <= x"ffaf07cd";
		wait for Clk_period;
		Addr <=  "0000111010101";
		Trees_din <= x"004b07cd";
		wait for Clk_period;
		Addr <=  "0000111010110";
		Trees_din <= x"400c5304";
		wait for Clk_period;
		Addr <=  "0000111010111";
		Trees_din <= x"ff6707cd";
		wait for Clk_period;
		Addr <=  "0000111011000";
		Trees_din <= x"001d07cd";
		wait for Clk_period;
		Addr <=  "0000111011001";
		Trees_din <= x"d7031d10";
		wait for Clk_period;
		Addr <=  "0000111011010";
		Trees_din <= x"01036508";
		wait for Clk_period;
		Addr <=  "0000111011011";
		Trees_din <= x"80026204";
		wait for Clk_period;
		Addr <=  "0000111011100";
		Trees_din <= x"ffe307cd";
		wait for Clk_period;
		Addr <=  "0000111011101";
		Trees_din <= x"00a007cd";
		wait for Clk_period;
		Addr <=  "0000111011110";
		Trees_din <= x"4d073b04";
		wait for Clk_period;
		Addr <=  "0000111011111";
		Trees_din <= x"ffa207cd";
		wait for Clk_period;
		Addr <=  "0000111100000";
		Trees_din <= x"fffe07cd";
		wait for Clk_period;
		Addr <=  "0000111100001";
		Trees_din <= x"36071f04";
		wait for Clk_period;
		Addr <=  "0000111100010";
		Trees_din <= x"ff7407cd";
		wait for Clk_period;
		Addr <=  "0000111100011";
		Trees_din <= x"6007f404";
		wait for Clk_period;
		Addr <=  "0000111100100";
		Trees_din <= x"004707cd";
		wait for Clk_period;
		Addr <=  "0000111100101";
		Trees_din <= x"ffa207cd";
		wait for Clk_period;
		Addr <=  "0000111100110";
		Trees_din <= x"4505d314";
		wait for Clk_period;
		Addr <=  "0000111100111";
		Trees_din <= x"4d040304";
		wait for Clk_period;
		Addr <=  "0000111101000";
		Trees_din <= x"ffae07cd";
		wait for Clk_period;
		Addr <=  "0000111101001";
		Trees_din <= x"42090d0c";
		wait for Clk_period;
		Addr <=  "0000111101010";
		Trees_din <= x"9b026f08";
		wait for Clk_period;
		Addr <=  "0000111101011";
		Trees_din <= x"3a019604";
		wait for Clk_period;
		Addr <=  "0000111101100";
		Trees_din <= x"00ba07cd";
		wait for Clk_period;
		Addr <=  "0000111101101";
		Trees_din <= x"003207cd";
		wait for Clk_period;
		Addr <=  "0000111101110";
		Trees_din <= x"001807cd";
		wait for Clk_period;
		Addr <=  "0000111101111";
		Trees_din <= x"fff607cd";
		wait for Clk_period;
		Addr <=  "0000111110000";
		Trees_din <= x"44030904";
		wait for Clk_period;
		Addr <=  "0000111110001";
		Trees_din <= x"002707cd";
		wait for Clk_period;
		Addr <=  "0000111110010";
		Trees_din <= x"ff8407cd";
		wait for Clk_period;
		Addr <=  "0000111110011";
		Trees_din <= x"1b074b28";
		wait for Clk_period;
		Addr <=  "0000111110100";
		Trees_din <= x"27067110";
		wait for Clk_period;
		Addr <=  "0000111110101";
		Trees_din <= x"97000104";
		wait for Clk_period;
		Addr <=  "0000111110110";
		Trees_din <= x"001a0849";
		wait for Clk_period;
		Addr <=  "0000111110111";
		Trees_din <= x"b7000104";
		wait for Clk_period;
		Addr <=  "0000111111000";
		Trees_din <= x"00060849";
		wait for Clk_period;
		Addr <=  "0000111111001";
		Trees_din <= x"3e0a8e04";
		wait for Clk_period;
		Addr <=  "0000111111010";
		Trees_din <= x"ff670849";
		wait for Clk_period;
		Addr <=  "0000111111011";
		Trees_din <= x"ffee0849";
		wait for Clk_period;
		Addr <=  "0000111111100";
		Trees_din <= x"16087c14";
		wait for Clk_period;
		Addr <=  "0000111111101";
		Trees_din <= x"1f05cb0c";
		wait for Clk_period;
		Addr <=  "0000111111110";
		Trees_din <= x"5e01e308";
		wait for Clk_period;
		Addr <=  "0000111111111";
		Trees_din <= x"01036504";
		wait for Clk_period;
		Addr <=  "0001000000000";
		Trees_din <= x"008e0849";
		wait for Clk_period;
		Addr <=  "0001000000001";
		Trees_din <= x"00010849";
		wait for Clk_period;
		Addr <=  "0001000000010";
		Trees_din <= x"ffba0849";
		wait for Clk_period;
		Addr <=  "0001000000011";
		Trees_din <= x"d9029c04";
		wait for Clk_period;
		Addr <=  "0001000000100";
		Trees_din <= x"fff10849";
		wait for Clk_period;
		Addr <=  "0001000000101";
		Trees_din <= x"ff930849";
		wait for Clk_period;
		Addr <=  "0001000000110";
		Trees_din <= x"ff790849";
		wait for Clk_period;
		Addr <=  "0001000000111";
		Trees_din <= x"45058210";
		wait for Clk_period;
		Addr <=  "0001000001000";
		Trees_din <= x"4d040304";
		wait for Clk_period;
		Addr <=  "0001000001001";
		Trees_din <= x"ffb70849";
		wait for Clk_period;
		Addr <=  "0001000001010";
		Trees_din <= x"42090d08";
		wait for Clk_period;
		Addr <=  "0001000001011";
		Trees_din <= x"3a019604";
		wait for Clk_period;
		Addr <=  "0001000001100";
		Trees_din <= x"00a70849";
		wait for Clk_period;
		Addr <=  "0001000001101";
		Trees_din <= x"00200849";
		wait for Clk_period;
		Addr <=  "0001000001110";
		Trees_din <= x"fffc0849";
		wait for Clk_period;
		Addr <=  "0001000001111";
		Trees_din <= x"270d9804";
		wait for Clk_period;
		Addr <=  "0001000010000";
		Trees_din <= x"ff880849";
		wait for Clk_period;
		Addr <=  "0001000010001";
		Trees_din <= x"00390849";
		wait for Clk_period;
		Addr <=  "0001000010010";
		Trees_din <= x"6b055718";
		wait for Clk_period;
		Addr <=  "0001000010011";
		Trees_din <= x"ba08eb0c";
		wait for Clk_period;
		Addr <=  "0001000010100";
		Trees_din <= x"1b087904";
		wait for Clk_period;
		Addr <=  "0001000010101";
		Trees_din <= x"ff6808c5";
		wait for Clk_period;
		Addr <=  "0001000010110";
		Trees_din <= x"7c006e04";
		wait for Clk_period;
		Addr <=  "0001000010111";
		Trees_din <= x"003f08c5";
		wait for Clk_period;
		Addr <=  "0001000011000";
		Trees_din <= x"ffb208c5";
		wait for Clk_period;
		Addr <=  "0001000011001";
		Trees_din <= x"8d02d604";
		wait for Clk_period;
		Addr <=  "0001000011010";
		Trees_din <= x"ff8908c5";
		wait for Clk_period;
		Addr <=  "0001000011011";
		Trees_din <= x"3b06e404";
		wait for Clk_period;
		Addr <=  "0001000011100";
		Trees_din <= x"001808c5";
		wait for Clk_period;
		Addr <=  "0001000011101";
		Trees_din <= x"007208c5";
		wait for Clk_period;
		Addr <=  "0001000011110";
		Trees_din <= x"1b035b10";
		wait for Clk_period;
		Addr <=  "0001000011111";
		Trees_din <= x"7e098908";
		wait for Clk_period;
		Addr <=  "0001000100000";
		Trees_din <= x"5205dd04";
		wait for Clk_period;
		Addr <=  "0001000100001";
		Trees_din <= x"ff7808c5";
		wait for Clk_period;
		Addr <=  "0001000100010";
		Trees_din <= x"fff208c5";
		wait for Clk_period;
		Addr <=  "0001000100011";
		Trees_din <= x"3401f704";
		wait for Clk_period;
		Addr <=  "0001000100100";
		Trees_din <= x"006d08c5";
		wait for Clk_period;
		Addr <=  "0001000100101";
		Trees_din <= x"ffa808c5";
		wait for Clk_period;
		Addr <=  "0001000100110";
		Trees_din <= x"c202110c";
		wait for Clk_period;
		Addr <=  "0001000100111";
		Trees_din <= x"8d014804";
		wait for Clk_period;
		Addr <=  "0001000101000";
		Trees_din <= x"000f08c5";
		wait for Clk_period;
		Addr <=  "0001000101001";
		Trees_din <= x"df04ac04";
		wait for Clk_period;
		Addr <=  "0001000101010";
		Trees_din <= x"003208c5";
		wait for Clk_period;
		Addr <=  "0001000101011";
		Trees_din <= x"00c708c5";
		wait for Clk_period;
		Addr <=  "0001000101100";
		Trees_din <= x"27062304";
		wait for Clk_period;
		Addr <=  "0001000101101";
		Trees_din <= x"ff8c08c5";
		wait for Clk_period;
		Addr <=  "0001000101110";
		Trees_din <= x"3201e704";
		wait for Clk_period;
		Addr <=  "0001000101111";
		Trees_din <= x"006f08c5";
		wait for Clk_period;
		Addr <=  "0001000110000";
		Trees_din <= x"fff508c5";
		wait for Clk_period;
		Addr <=  "0001000110001";
		Trees_din <= x"6b055710";
		wait for Clk_period;
		Addr <=  "0001000110010";
		Trees_din <= x"ba08eb08";
		wait for Clk_period;
		Addr <=  "0001000110011";
		Trees_din <= x"d1002004";
		wait for Clk_period;
		Addr <=  "0001000110100";
		Trees_din <= x"fffd0929";
		wait for Clk_period;
		Addr <=  "0001000110101";
		Trees_din <= x"ff690929";
		wait for Clk_period;
		Addr <=  "0001000110110";
		Trees_din <= x"8d02d604";
		wait for Clk_period;
		Addr <=  "0001000110111";
		Trees_din <= x"ff900929";
		wait for Clk_period;
		Addr <=  "0001000111000";
		Trees_din <= x"00570929";
		wait for Clk_period;
		Addr <=  "0001000111001";
		Trees_din <= x"34023414";
		wait for Clk_period;
		Addr <=  "0001000111010";
		Trees_din <= x"38058510";
		wait for Clk_period;
		Addr <=  "0001000111011";
		Trees_din <= x"c201e608";
		wait for Clk_period;
		Addr <=  "0001000111100";
		Trees_din <= x"17018304";
		wait for Clk_period;
		Addr <=  "0001000111101";
		Trees_din <= x"00c00929";
		wait for Clk_period;
		Addr <=  "0001000111110";
		Trees_din <= x"002c0929";
		wait for Clk_period;
		Addr <=  "0001000111111";
		Trees_din <= x"6b0c7104";
		wait for Clk_period;
		Addr <=  "0001001000000";
		Trees_din <= x"ffcf0929";
		wait for Clk_period;
		Addr <=  "0001001000001";
		Trees_din <= x"00500929";
		wait for Clk_period;
		Addr <=  "0001001000010";
		Trees_din <= x"ffa70929";
		wait for Clk_period;
		Addr <=  "0001001000011";
		Trees_din <= x"360afc08";
		wait for Clk_period;
		Addr <=  "0001001000100";
		Trees_din <= x"58059304";
		wait for Clk_period;
		Addr <=  "0001001000101";
		Trees_din <= x"ff810929";
		wait for Clk_period;
		Addr <=  "0001001000110";
		Trees_din <= x"00120929";
		wait for Clk_period;
		Addr <=  "0001001000111";
		Trees_din <= x"3504d404";
		wait for Clk_period;
		Addr <=  "0001001001000";
		Trees_din <= x"fffe0929";
		wait for Clk_period;
		Addr <=  "0001001001001";
		Trees_din <= x"00460929";
		wait for Clk_period;
		Addr <=  "0001001001010";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0001001001011";
		Trees_din <= x"6b055714";
		wait for Clk_period;
		Addr <=  "0001001001100";
		Trees_din <= x"02067b08";
		wait for Clk_period;
		Addr <=  "0001001001101";
		Trees_din <= x"dc0d3304";
		wait for Clk_period;
		Addr <=  "0001001001110";
		Trees_din <= x"ff6b0989";
		wait for Clk_period;
		Addr <=  "0001001001111";
		Trees_din <= x"ffd40989";
		wait for Clk_period;
		Addr <=  "0001001010000";
		Trees_din <= x"13031f08";
		wait for Clk_period;
		Addr <=  "0001001010001";
		Trees_din <= x"1b051e04";
		wait for Clk_period;
		Addr <=  "0001001010010";
		Trees_din <= x"ffdf0989";
		wait for Clk_period;
		Addr <=  "0001001010011";
		Trees_din <= x"006c0989";
		wait for Clk_period;
		Addr <=  "0001001010100";
		Trees_din <= x"ff8b0989";
		wait for Clk_period;
		Addr <=  "0001001010101";
		Trees_din <= x"1b035b0c";
		wait for Clk_period;
		Addr <=  "0001001010110";
		Trees_din <= x"7e098908";
		wait for Clk_period;
		Addr <=  "0001001010111";
		Trees_din <= x"52046004";
		wait for Clk_period;
		Addr <=  "0001001011000";
		Trees_din <= x"ff810989";
		wait for Clk_period;
		Addr <=  "0001001011001";
		Trees_din <= x"ffe50989";
		wait for Clk_period;
		Addr <=  "0001001011010";
		Trees_din <= x"000e0989";
		wait for Clk_period;
		Addr <=  "0001001011011";
		Trees_din <= x"3804020c";
		wait for Clk_period;
		Addr <=  "0001001011100";
		Trees_din <= x"0d029408";
		wait for Clk_period;
		Addr <=  "0001001011101";
		Trees_din <= x"1c02a604";
		wait for Clk_period;
		Addr <=  "0001001011110";
		Trees_din <= x"00290989";
		wait for Clk_period;
		Addr <=  "0001001011111";
		Trees_din <= x"00a80989";
		wait for Clk_period;
		Addr <=  "0001001100000";
		Trees_din <= x"fff10989";
		wait for Clk_period;
		Addr <=  "0001001100001";
		Trees_din <= x"ffb40989";
		wait for Clk_period;
		Addr <=  "0001001100010";
		Trees_din <= x"6b055710";
		wait for Clk_period;
		Addr <=  "0001001100011";
		Trees_din <= x"1c073008";
		wait for Clk_period;
		Addr <=  "0001001100100";
		Trees_din <= x"360afc04";
		wait for Clk_period;
		Addr <=  "0001001100101";
		Trees_din <= x"ff6f09e5";
		wait for Clk_period;
		Addr <=  "0001001100110";
		Trees_din <= x"000f09e5";
		wait for Clk_period;
		Addr <=  "0001001100111";
		Trees_din <= x"fd02e204";
		wait for Clk_period;
		Addr <=  "0001001101000";
		Trees_din <= x"ffb109e5";
		wait for Clk_period;
		Addr <=  "0001001101001";
		Trees_din <= x"005609e5";
		wait for Clk_period;
		Addr <=  "0001001101010";
		Trees_din <= x"34023410";
		wait for Clk_period;
		Addr <=  "0001001101011";
		Trees_din <= x"1504230c";
		wait for Clk_period;
		Addr <=  "0001001101100";
		Trees_din <= x"c201e608";
		wait for Clk_period;
		Addr <=  "0001001101101";
		Trees_din <= x"5c019804";
		wait for Clk_period;
		Addr <=  "0001001101110";
		Trees_din <= x"002909e5";
		wait for Clk_period;
		Addr <=  "0001001101111";
		Trees_din <= x"00ae09e5";
		wait for Clk_period;
		Addr <=  "0001001110000";
		Trees_din <= x"001509e5";
		wait for Clk_period;
		Addr <=  "0001001110001";
		Trees_din <= x"ffc809e5";
		wait for Clk_period;
		Addr <=  "0001001110010";
		Trees_din <= x"7a072d08";
		wait for Clk_period;
		Addr <=  "0001001110011";
		Trees_din <= x"58050e04";
		wait for Clk_period;
		Addr <=  "0001001110100";
		Trees_din <= x"ff8209e5";
		wait for Clk_period;
		Addr <=  "0001001110101";
		Trees_din <= x"000809e5";
		wait for Clk_period;
		Addr <=  "0001001110110";
		Trees_din <= x"1b06ce04";
		wait for Clk_period;
		Addr <=  "0001001110111";
		Trees_din <= x"ffdd09e5";
		wait for Clk_period;
		Addr <=  "0001001111000";
		Trees_din <= x"004909e5";
		wait for Clk_period;
		Addr <=  "0001001111001";
		Trees_din <= x"7504ce0c";
		wait for Clk_period;
		Addr <=  "0001001111010";
		Trees_din <= x"720a4708";
		wait for Clk_period;
		Addr <=  "0001001111011";
		Trees_din <= x"27074404";
		wait for Clk_period;
		Addr <=  "0001001111100";
		Trees_din <= x"ff710a31";
		wait for Clk_period;
		Addr <=  "0001001111101";
		Trees_din <= x"fff50a31";
		wait for Clk_period;
		Addr <=  "0001001111110";
		Trees_din <= x"00300a31";
		wait for Clk_period;
		Addr <=  "0001001111111";
		Trees_din <= x"1c02c00c";
		wait for Clk_period;
		Addr <=  "0001010000000";
		Trees_din <= x"0400bc04";
		wait for Clk_period;
		Addr <=  "0001010000001";
		Trees_din <= x"000c0a31";
		wait for Clk_period;
		Addr <=  "0001010000010";
		Trees_din <= x"7b04ef04";
		wait for Clk_period;
		Addr <=  "0001010000011";
		Trees_din <= x"ff880a31";
		wait for Clk_period;
		Addr <=  "0001010000100";
		Trees_din <= x"ffe50a31";
		wait for Clk_period;
		Addr <=  "0001010000101";
		Trees_din <= x"b5025d0c";
		wait for Clk_period;
		Addr <=  "0001010000110";
		Trees_din <= x"01053a08";
		wait for Clk_period;
		Addr <=  "0001010000111";
		Trees_din <= x"17019904";
		wait for Clk_period;
		Addr <=  "0001010001000";
		Trees_din <= x"00a30a31";
		wait for Clk_period;
		Addr <=  "0001010001001";
		Trees_din <= x"002a0a31";
		wait for Clk_period;
		Addr <=  "0001010001010";
		Trees_din <= x"fff30a31";
		wait for Clk_period;
		Addr <=  "0001010001011";
		Trees_din <= x"ffaf0a31";
		wait for Clk_period;
		Addr <=  "0001010001100";
		Trees_din <= x"6b055714";
		wait for Clk_period;
		Addr <=  "0001010001101";
		Trees_din <= x"02067b08";
		wait for Clk_period;
		Addr <=  "0001010001110";
		Trees_din <= x"36071f04";
		wait for Clk_period;
		Addr <=  "0001010001111";
		Trees_din <= x"ff700a85";
		wait for Clk_period;
		Addr <=  "0001010010000";
		Trees_din <= x"ffd50a85";
		wait for Clk_period;
		Addr <=  "0001010010001";
		Trees_din <= x"01020c08";
		wait for Clk_period;
		Addr <=  "0001010010010";
		Trees_din <= x"1c073004";
		wait for Clk_period;
		Addr <=  "0001010010011";
		Trees_din <= x"00080a85";
		wait for Clk_period;
		Addr <=  "0001010010100";
		Trees_din <= x"00540a85";
		wait for Clk_period;
		Addr <=  "0001010010101";
		Trees_din <= x"ffa00a85";
		wait for Clk_period;
		Addr <=  "0001010010110";
		Trees_din <= x"1b035b08";
		wait for Clk_period;
		Addr <=  "0001010010111";
		Trees_din <= x"7e098904";
		wait for Clk_period;
		Addr <=  "0001010011000";
		Trees_din <= x"ff9d0a85";
		wait for Clk_period;
		Addr <=  "0001010011001";
		Trees_din <= x"000d0a85";
		wait for Clk_period;
		Addr <=  "0001010011010";
		Trees_din <= x"3801ea08";
		wait for Clk_period;
		Addr <=  "0001010011011";
		Trees_din <= x"0d01d704";
		wait for Clk_period;
		Addr <=  "0001010011100";
		Trees_din <= x"00900a85";
		wait for Clk_period;
		Addr <=  "0001010011101";
		Trees_din <= x"00100a85";
		wait for Clk_period;
		Addr <=  "0001010011110";
		Trees_din <= x"c10b8704";
		wait for Clk_period;
		Addr <=  "0001010011111";
		Trees_din <= x"ffba0a85";
		wait for Clk_period;
		Addr <=  "0001010100000";
		Trees_din <= x"00250a85";
		wait for Clk_period;
		Addr <=  "0001010100001";
		Trees_din <= x"6b055710";
		wait for Clk_period;
		Addr <=  "0001010100010";
		Trees_din <= x"7d00ad08";
		wait for Clk_period;
		Addr <=  "0001010100011";
		Trees_din <= x"8d02f304";
		wait for Clk_period;
		Addr <=  "0001010100100";
		Trees_din <= x"ffac0ad1";
		wait for Clk_period;
		Addr <=  "0001010100101";
		Trees_din <= x"002f0ad1";
		wait for Clk_period;
		Addr <=  "0001010100110";
		Trees_din <= x"36070204";
		wait for Clk_period;
		Addr <=  "0001010100111";
		Trees_din <= x"ff730ad1";
		wait for Clk_period;
		Addr <=  "0001010101000";
		Trees_din <= x"ffda0ad1";
		wait for Clk_period;
		Addr <=  "0001010101001";
		Trees_din <= x"df04e20c";
		wait for Clk_period;
		Addr <=  "0001010101010";
		Trees_din <= x"35054f04";
		wait for Clk_period;
		Addr <=  "0001010101011";
		Trees_din <= x"ff9a0ad1";
		wait for Clk_period;
		Addr <=  "0001010101100";
		Trees_din <= x"4f021504";
		wait for Clk_period;
		Addr <=  "0001010101101";
		Trees_din <= x"ffd10ad1";
		wait for Clk_period;
		Addr <=  "0001010101110";
		Trees_din <= x"00320ad1";
		wait for Clk_period;
		Addr <=  "0001010101111";
		Trees_din <= x"3404b808";
		wait for Clk_period;
		Addr <=  "0001010110000";
		Trees_din <= x"01031804";
		wait for Clk_period;
		Addr <=  "0001010110001";
		Trees_din <= x"00850ad1";
		wait for Clk_period;
		Addr <=  "0001010110010";
		Trees_din <= x"001b0ad1";
		wait for Clk_period;
		Addr <=  "0001010110011";
		Trees_din <= x"ffd90ad1";
		wait for Clk_period;
		Addr <=  "0001010110100";
		Trees_din <= x"1b03870c";
		wait for Clk_period;
		Addr <=  "0001010110101";
		Trees_din <= x"98080704";
		wait for Clk_period;
		Addr <=  "0001010110110";
		Trees_din <= x"ff7d0b15";
		wait for Clk_period;
		Addr <=  "0001010110111";
		Trees_din <= x"34026604";
		wait for Clk_period;
		Addr <=  "0001010111000";
		Trees_din <= x"00370b15";
		wait for Clk_period;
		Addr <=  "0001010111001";
		Trees_din <= x"ffb70b15";
		wait for Clk_period;
		Addr <=  "0001010111010";
		Trees_din <= x"7505860c";
		wait for Clk_period;
		Addr <=  "0001010111011";
		Trees_din <= x"3801f708";
		wait for Clk_period;
		Addr <=  "0001010111100";
		Trees_din <= x"de00fb04";
		wait for Clk_period;
		Addr <=  "0001010111101";
		Trees_din <= x"003d0b15";
		wait for Clk_period;
		Addr <=  "0001010111110";
		Trees_din <= x"ffda0b15";
		wait for Clk_period;
		Addr <=  "0001010111111";
		Trees_din <= x"ff990b15";
		wait for Clk_period;
		Addr <=  "0001011000000";
		Trees_din <= x"45058208";
		wait for Clk_period;
		Addr <=  "0001011000001";
		Trees_din <= x"a4041204";
		wait for Clk_period;
		Addr <=  "0001011000010";
		Trees_din <= x"00800b15";
		wait for Clk_period;
		Addr <=  "0001011000011";
		Trees_din <= x"001d0b15";
		wait for Clk_period;
		Addr <=  "0001011000100";
		Trees_din <= x"ffe00b15";
		wait for Clk_period;
		Addr <=  "0001011000101";
		Trees_din <= x"36070214";
		wait for Clk_period;
		Addr <=  "0001011000110";
		Trees_din <= x"9b007408";
		wait for Clk_period;
		Addr <=  "0001011000111";
		Trees_din <= x"1e06cf04";
		wait for Clk_period;
		Addr <=  "0001011001000";
		Trees_din <= x"ffd90b51";
		wait for Clk_period;
		Addr <=  "0001011001001";
		Trees_din <= x"004f0b51";
		wait for Clk_period;
		Addr <=  "0001011001010";
		Trees_din <= x"1c073008";
		wait for Clk_period;
		Addr <=  "0001011001011";
		Trees_din <= x"6b094104";
		wait for Clk_period;
		Addr <=  "0001011001100";
		Trees_din <= x"ff780b51";
		wait for Clk_period;
		Addr <=  "0001011001101";
		Trees_din <= x"ffda0b51";
		wait for Clk_period;
		Addr <=  "0001011001110";
		Trees_din <= x"00180b51";
		wait for Clk_period;
		Addr <=  "0001011001111";
		Trees_din <= x"3404b808";
		wait for Clk_period;
		Addr <=  "0001011010000";
		Trees_din <= x"2103de04";
		wait for Clk_period;
		Addr <=  "0001011010001";
		Trees_din <= x"ffff0b51";
		wait for Clk_period;
		Addr <=  "0001011010010";
		Trees_din <= x"005f0b51";
		wait for Clk_period;
		Addr <=  "0001011010011";
		Trees_din <= x"ffca0b51";
		wait for Clk_period;
		Addr <=  "0001011010100";
		Trees_din <= x"1b03870c";
		wait for Clk_period;
		Addr <=  "0001011010101";
		Trees_din <= x"94079504";
		wait for Clk_period;
		Addr <=  "0001011010110";
		Trees_din <= x"ff7f0b8d";
		wait for Clk_period;
		Addr <=  "0001011010111";
		Trees_din <= x"18015c04";
		wait for Clk_period;
		Addr <=  "0001011011000";
		Trees_din <= x"ffb40b8d";
		wait for Clk_period;
		Addr <=  "0001011011001";
		Trees_din <= x"00190b8d";
		wait for Clk_period;
		Addr <=  "0001011011010";
		Trees_din <= x"01021d0c";
		wait for Clk_period;
		Addr <=  "0001011011011";
		Trees_din <= x"29038308";
		wait for Clk_period;
		Addr <=  "0001011011100";
		Trees_din <= x"75048204";
		wait for Clk_period;
		Addr <=  "0001011011101";
		Trees_din <= x"001b0b8d";
		wait for Clk_period;
		Addr <=  "0001011011110";
		Trees_din <= x"00770b8d";
		wait for Clk_period;
		Addr <=  "0001011011111";
		Trees_din <= x"ffe70b8d";
		wait for Clk_period;
		Addr <=  "0001011100000";
		Trees_din <= x"2107e304";
		wait for Clk_period;
		Addr <=  "0001011100001";
		Trees_din <= x"ffa10b8d";
		wait for Clk_period;
		Addr <=  "0001011100010";
		Trees_din <= x"001e0b8d";
		wait for Clk_period;
		Addr <=  "0001011100011";
		Trees_din <= x"3801f70c";
		wait for Clk_period;
		Addr <=  "0001011100100";
		Trees_din <= x"b5025d08";
		wait for Clk_period;
		Addr <=  "0001011100101";
		Trees_din <= x"01036504";
		wait for Clk_period;
		Addr <=  "0001011100110";
		Trees_din <= x"00680bb1";
		wait for Clk_period;
		Addr <=  "0001011100111";
		Trees_din <= x"ffea0bb1";
		wait for Clk_period;
		Addr <=  "0001011101000";
		Trees_din <= x"ffa60bb1";
		wait for Clk_period;
		Addr <=  "0001011101001";
		Trees_din <= x"c10a0004";
		wait for Clk_period;
		Addr <=  "0001011101010";
		Trees_din <= x"ff870bb1";
		wait for Clk_period;
		Addr <=  "0001011101011";
		Trees_din <= x"00040bb1";
		wait for Clk_period;
		Addr <=  "0001011101100";
		Trees_din <= x"1b035b08";
		wait for Clk_period;
		Addr <=  "0001011101101";
		Trees_din <= x"36070204";
		wait for Clk_period;
		Addr <=  "0001011101110";
		Trees_din <= x"ff910bdd";
		wait for Clk_period;
		Addr <=  "0001011101111";
		Trees_din <= x"00010bdd";
		wait for Clk_period;
		Addr <=  "0001011110000";
		Trees_din <= x"3802d30c";
		wait for Clk_period;
		Addr <=  "0001011110001";
		Trees_din <= x"13038a08";
		wait for Clk_period;
		Addr <=  "0001011110010";
		Trees_din <= x"17016204";
		wait for Clk_period;
		Addr <=  "0001011110011";
		Trees_din <= x"006b0bdd";
		wait for Clk_period;
		Addr <=  "0001011110100";
		Trees_din <= x"00080bdd";
		wait for Clk_period;
		Addr <=  "0001011110101";
		Trees_din <= x"ffe50bdd";
		wait for Clk_period;
		Addr <=  "0001011110110";
		Trees_din <= x"ffc00bdd";
		wait for Clk_period;
		Addr <=  "0001011110111";
		Trees_din <= x"6b055708";
		wait for Clk_period;
		Addr <=  "0001011111000";
		Trees_din <= x"11075004";
		wait for Clk_period;
		Addr <=  "0001011111001";
		Trees_din <= x"ff900c01";
		wait for Clk_period;
		Addr <=  "0001011111010";
		Trees_din <= x"00040c01";
		wait for Clk_period;
		Addr <=  "0001011111011";
		Trees_din <= x"3404b808";
		wait for Clk_period;
		Addr <=  "0001011111100";
		Trees_din <= x"1c02c004";
		wait for Clk_period;
		Addr <=  "0001011111101";
		Trees_din <= x"fffb0c01";
		wait for Clk_period;
		Addr <=  "0001011111110";
		Trees_din <= x"00540c01";
		wait for Clk_period;
		Addr <=  "0001011111111";
		Trees_din <= x"ffc60c01";
		wait for Clk_period;
		Addr <=  "0001100000000";
		Trees_din <= x"3801f70c";
		wait for Clk_period;
		Addr <=  "0001100000001";
		Trees_din <= x"17016208";
		wait for Clk_period;
		Addr <=  "0001100000010";
		Trees_din <= x"8d02ed04";
		wait for Clk_period;
		Addr <=  "0001100000011";
		Trees_din <= x"00090c25";
		wait for Clk_period;
		Addr <=  "0001100000100";
		Trees_din <= x"00560c25";
		wait for Clk_period;
		Addr <=  "0001100000101";
		Trees_din <= x"ffdd0c25";
		wait for Clk_period;
		Addr <=  "0001100000110";
		Trees_din <= x"270a8204";
		wait for Clk_period;
		Addr <=  "0001100000111";
		Trees_din <= x"ff9a0c25";
		wait for Clk_period;
		Addr <=  "0001100001000";
		Trees_din <= x"00120c25";
		wait for Clk_period;
		Addr <=  "0001100001001";
		Trees_din <= x"1b035b08";
		wait for Clk_period;
		Addr <=  "0001100001010";
		Trees_din <= x"a406f004";
		wait for Clk_period;
		Addr <=  "0001100001011";
		Trees_din <= x"ff9b0c49";
		wait for Clk_period;
		Addr <=  "0001100001100";
		Trees_din <= x"00000c49";
		wait for Clk_period;
		Addr <=  "0001100001101";
		Trees_din <= x"3802d308";
		wait for Clk_period;
		Addr <=  "0001100001110";
		Trees_din <= x"a4047704";
		wait for Clk_period;
		Addr <=  "0001100001111";
		Trees_din <= x"004d0c49";
		wait for Clk_period;
		Addr <=  "0001100010000";
		Trees_din <= x"fff60c49";
		wait for Clk_period;
		Addr <=  "0001100010001";
		Trees_din <= x"ffd00c49";
		wait for Clk_period;
		Addr <=  "0001100010010";
		Trees_din <= x"3b045808";
		wait for Clk_period;
		Addr <=  "0001100010011";
		Trees_din <= x"36071f04";
		wait for Clk_period;
		Addr <=  "0001100010100";
		Trees_din <= x"ffa10c65";
		wait for Clk_period;
		Addr <=  "0001100010101";
		Trees_din <= x"000b0c65";
		wait for Clk_period;
		Addr <=  "0001100010110";
		Trees_din <= x"fa024b04";
		wait for Clk_period;
		Addr <=  "0001100010111";
		Trees_din <= x"004a0c65";
		wait for Clk_period;
		Addr <=  "0001100011000";
		Trees_din <= x"ffdf0c65";
		wait for Clk_period;
		Addr <=  "0001100011001";
		Trees_din <= x"11042e08";
		wait for Clk_period;
		Addr <=  "0001100011010";
		Trees_din <= x"21054504";
		wait for Clk_period;
		Addr <=  "0001100011011";
		Trees_din <= x"ffa30c89";
		wait for Clk_period;
		Addr <=  "0001100011100";
		Trees_din <= x"ffee0c89";
		wait for Clk_period;
		Addr <=  "0001100011101";
		Trees_din <= x"45051308";
		wait for Clk_period;
		Addr <=  "0001100011110";
		Trees_din <= x"01021d04";
		wait for Clk_period;
		Addr <=  "0001100011111";
		Trees_din <= x"004e0c89";
		wait for Clk_period;
		Addr <=  "0001100100000";
		Trees_din <= x"fff90c89";
		wait for Clk_period;
		Addr <=  "0001100100001";
		Trees_din <= x"ffd00c89";
		wait for Clk_period;
		Addr <=  "0001100100010";
		Trees_din <= x"1b035b08";
		wait for Clk_period;
		Addr <=  "0001100100011";
		Trees_din <= x"27080204";
		wait for Clk_period;
		Addr <=  "0001100100100";
		Trees_din <= x"ffa30cad";
		wait for Clk_period;
		Addr <=  "0001100100101";
		Trees_din <= x"fff90cad";
		wait for Clk_period;
		Addr <=  "0001100100110";
		Trees_din <= x"13038a08";
		wait for Clk_period;
		Addr <=  "0001100100111";
		Trees_din <= x"3a012804";
		wait for Clk_period;
		Addr <=  "0001100101000";
		Trees_din <= x"00470cad";
		wait for Clk_period;
		Addr <=  "0001100101001";
		Trees_din <= x"00080cad";
		wait for Clk_period;
		Addr <=  "0001100101010";
		Trees_din <= x"ffe00cad";
		wait for Clk_period;
		Addr <=  "0001100101011";
		Trees_din <= x"01021d08";
		wait for Clk_period;
		Addr <=  "0001100101100";
		Trees_din <= x"cf020404";
		wait for Clk_period;
		Addr <=  "0001100101101";
		Trees_din <= x"00400cc9";
		wait for Clk_period;
		Addr <=  "0001100101110";
		Trees_din <= x"ffe30cc9";
		wait for Clk_period;
		Addr <=  "0001100101111";
		Trees_din <= x"27085d04";
		wait for Clk_period;
		Addr <=  "0001100110000";
		Trees_din <= x"ffa80cc9";
		wait for Clk_period;
		Addr <=  "0001100110001";
		Trees_din <= x"000a0cc9";
		wait for Clk_period;
		Addr <=  "0001100110010";
		Trees_din <= x"3605f808";
		wait for Clk_period;
		Addr <=  "0001100110011";
		Trees_din <= x"35054f04";
		wait for Clk_period;
		Addr <=  "0001100110100";
		Trees_din <= x"ffaf0ce5";
		wait for Clk_period;
		Addr <=  "0001100110101";
		Trees_din <= x"00090ce5";
		wait for Clk_period;
		Addr <=  "0001100110110";
		Trees_din <= x"1c042d04";
		wait for Clk_period;
		Addr <=  "0001100110111";
		Trees_din <= x"fffb0ce5";
		wait for Clk_period;
		Addr <=  "0001100111000";
		Trees_din <= x"00370ce5";
		wait for Clk_period;
		Addr <=  "0001100111001";
		Trees_din <= x"1c02c008";
		wait for Clk_period;
		Addr <=  "0001100111010";
		Trees_din <= x"68028b04";
		wait for Clk_period;
		Addr <=  "0001100111011";
		Trees_din <= x"ffb20d01";
		wait for Clk_period;
		Addr <=  "0001100111100";
		Trees_din <= x"fffa0d01";
		wait for Clk_period;
		Addr <=  "0001100111101";
		Trees_din <= x"75050b04";
		wait for Clk_period;
		Addr <=  "0001100111110";
		Trees_din <= x"ffe00d01";
		wait for Clk_period;
		Addr <=  "0001100111111";
		Trees_din <= x"003b0d01";
		wait for Clk_period;
		Addr <=  "0001101000000";
		Trees_din <= x"01021d08";
		wait for Clk_period;
		Addr <=  "0001101000001";
		Trees_din <= x"cf01e504";
		wait for Clk_period;
		Addr <=  "0001101000010";
		Trees_din <= x"003a0d1d";
		wait for Clk_period;
		Addr <=  "0001101000011";
		Trees_din <= x"ffec0d1d";
		wait for Clk_period;
		Addr <=  "0001101000100";
		Trees_din <= x"fd09aa04";
		wait for Clk_period;
		Addr <=  "0001101000101";
		Trees_din <= x"ffb10d1d";
		wait for Clk_period;
		Addr <=  "0001101000110";
		Trees_din <= x"00050d1d";
		wait for Clk_period;
		Addr <=  "0001101000111";
		Trees_din <= x"3402da08";
		wait for Clk_period;
		Addr <=  "0001101001000";
		Trees_din <= x"17018304";
		wait for Clk_period;
		Addr <=  "0001101001001";
		Trees_din <= x"00350d31";
		wait for Clk_period;
		Addr <=  "0001101001010";
		Trees_din <= x"ffe80d31";
		wait for Clk_period;
		Addr <=  "0001101001011";
		Trees_din <= x"ffcb0d31";
		wait for Clk_period;
		Addr <=  "0001101001100";
		Trees_din <= x"1b035b04";
		wait for Clk_period;
		Addr <=  "0001101001101";
		Trees_din <= x"ffcc0d45";
		wait for Clk_period;
		Addr <=  "0001101001110";
		Trees_din <= x"21049104";
		wait for Clk_period;
		Addr <=  "0001101001111";
		Trees_din <= x"ffed0d45";
		wait for Clk_period;
		Addr <=  "0001101010000";
		Trees_din <= x"00320d45";
		wait for Clk_period;
		Addr <=  "0001101010001";
		Trees_din <= x"01021d08";
		wait for Clk_period;
		Addr <=  "0001101010010";
		Trees_din <= x"cf014f04";
		wait for Clk_period;
		Addr <=  "0001101010011";
		Trees_din <= x"00370d59";
		wait for Clk_period;
		Addr <=  "0001101010100";
		Trees_din <= x"fff80d59";
		wait for Clk_period;
		Addr <=  "0001101010101";
		Trees_din <= x"ffd20d59";
		wait for Clk_period;
		Addr <=  "0001101010110";
		Trees_din <= x"7d011008";
		wait for Clk_period;
		Addr <=  "0001101010111";
		Trees_din <= x"1c043704";
		wait for Clk_period;
		Addr <=  "0001101011000";
		Trees_din <= x"fff70d6d";
		wait for Clk_period;
		Addr <=  "0001101011001";
		Trees_din <= x"00300d6d";
		wait for Clk_period;
		Addr <=  "0001101011010";
		Trees_din <= x"ffd20d6d";
		wait for Clk_period;
		Addr <=  "0001101011011";
		Trees_din <= x"3801f708";
		wait for Clk_period;
		Addr <=  "0001101011100";
		Trees_din <= x"4702c704";
		wait for Clk_period;
		Addr <=  "0001101011101";
		Trees_din <= x"002c0d81";
		wait for Clk_period;
		Addr <=  "0001101011110";
		Trees_din <= x"00000d81";
		wait for Clk_period;
		Addr <=  "0001101011111";
		Trees_din <= x"ffd70d81";
		wait for Clk_period;
		Addr <=  "0001101100000";
		Trees_din <= x"3402da08";
		wait for Clk_period;
		Addr <=  "0001101100001";
		Trees_din <= x"df058804";
		wait for Clk_period;
		Addr <=  "0001101100010";
		Trees_din <= x"fff70d95";
		wait for Clk_period;
		Addr <=  "0001101100011";
		Trees_din <= x"00300d95";
		wait for Clk_period;
		Addr <=  "0001101100100";
		Trees_din <= x"ffd40d95";
		wait for Clk_period;
		Addr <=  "0001101100101";
		Trees_din <= x"3605f804";
		wait for Clk_period;
		Addr <=  "0001101100110";
		Trees_din <= x"ffdb0da1";
		wait for Clk_period;
		Addr <=  "0001101100111";
		Trees_din <= x"001f0da1";
		wait for Clk_period;
		Addr <=  "0001101101000";
		Trees_din <= x"0000000f";
		wait for Clk_period;

        -- Class  6
        -----------
		Addr <=  "0000000000000";
		Trees_din <= x"1a0da620";
		wait for Clk_period;
		Addr <=  "0000000000001";
		Trees_din <= x"17136018";
		wait for Clk_period;
		Addr <=  "0000000000010";
		Trees_din <= x"71116a14";
		wait for Clk_period;
		Addr <=  "0000000000011";
		Trees_din <= x"190e0010";
		wait for Clk_period;
		Addr <=  "0000000000100";
		Trees_din <= x"1a096808";
		wait for Clk_period;
		Addr <=  "0000000000101";
		Trees_din <= x"770e7104";
		wait for Clk_period;
		Addr <=  "0000000000110";
		Trees_din <= x"ff4d004d";
		wait for Clk_period;
		Addr <=  "0000000000111";
		Trees_din <= x"ffb5004d";
		wait for Clk_period;
		Addr <=  "0000000001000";
		Trees_din <= x"db010104";
		wait for Clk_period;
		Addr <=  "0000000001001";
		Trees_din <= x"0164004d";
		wait for Clk_period;
		Addr <=  "0000000001010";
		Trees_din <= x"ff5c004d";
		wait for Clk_period;
		Addr <=  "0000000001011";
		Trees_din <= x"00a4004d";
		wait for Clk_period;
		Addr <=  "0000000001100";
		Trees_din <= x"00e2004d";
		wait for Clk_period;
		Addr <=  "0000000001101";
		Trees_din <= x"1a02a104";
		wait for Clk_period;
		Addr <=  "0000000001110";
		Trees_din <= x"ff8f004d";
		wait for Clk_period;
		Addr <=  "0000000001111";
		Trees_din <= x"02e4004d";
		wait for Clk_period;
		Addr <=  "0000000010000";
		Trees_din <= x"52010004";
		wait for Clk_period;
		Addr <=  "0000000010001";
		Trees_din <= x"fff1004d";
		wait for Clk_period;
		Addr <=  "0000000010010";
		Trees_din <= x"0403004d";
		wait for Clk_period;
		Addr <=  "0000000010011";
		Trees_din <= x"1a0acd24";
		wait for Clk_period;
		Addr <=  "0000000010100";
		Trees_din <= x"1713601c";
		wait for Clk_period;
		Addr <=  "0000000010101";
		Trees_din <= x"190e0014";
		wait for Clk_period;
		Addr <=  "0000000010110";
		Trees_din <= x"71116a10";
		wait for Clk_period;
		Addr <=  "0000000010111";
		Trees_din <= x"1a096808";
		wait for Clk_period;
		Addr <=  "0000000011000";
		Trees_din <= x"770e7104";
		wait for Clk_period;
		Addr <=  "0000000011001";
		Trees_din <= x"ff5400b9";
		wait for Clk_period;
		Addr <=  "0000000011010";
		Trees_din <= x"ffc200b9";
		wait for Clk_period;
		Addr <=  "0000000011011";
		Trees_din <= x"1b007704";
		wait for Clk_period;
		Addr <=  "0000000011100";
		Trees_din <= x"00cf00b9";
		wait for Clk_period;
		Addr <=  "0000000011101";
		Trees_din <= x"ff6d00b9";
		wait for Clk_period;
		Addr <=  "0000000011110";
		Trees_din <= x"001600b9";
		wait for Clk_period;
		Addr <=  "0000000011111";
		Trees_din <= x"1705e104";
		wait for Clk_period;
		Addr <=  "0000000100000";
		Trees_din <= x"ff9d00b9";
		wait for Clk_period;
		Addr <=  "0000000100001";
		Trees_din <= x"015d00b9";
		wait for Clk_period;
		Addr <=  "0000000100010";
		Trees_din <= x"1a02a104";
		wait for Clk_period;
		Addr <=  "0000000100011";
		Trees_din <= x"ff9b00b9";
		wait for Clk_period;
		Addr <=  "0000000100100";
		Trees_din <= x"019500b9";
		wait for Clk_period;
		Addr <=  "0000000100101";
		Trees_din <= x"17087b08";
		wait for Clk_period;
		Addr <=  "0000000100110";
		Trees_din <= x"06017604";
		wait for Clk_period;
		Addr <=  "0000000100111";
		Trees_din <= x"00b200b9";
		wait for Clk_period;
		Addr <=  "0000000101000";
		Trees_din <= x"ff7000b9";
		wait for Clk_period;
		Addr <=  "0000000101001";
		Trees_din <= x"43055104";
		wait for Clk_period;
		Addr <=  "0000000101010";
		Trees_din <= x"001b00b9";
		wait for Clk_period;
		Addr <=  "0000000101011";
		Trees_din <= x"0f073b04";
		wait for Clk_period;
		Addr <=  "0000000101100";
		Trees_din <= x"01c800b9";
		wait for Clk_period;
		Addr <=  "0000000101101";
		Trees_din <= x"009300b9";
		wait for Clk_period;
		Addr <=  "0000000101110";
		Trees_din <= x"1a0acd1c";
		wait for Clk_period;
		Addr <=  "0000000101111";
		Trees_din <= x"170de110";
		wait for Clk_period;
		Addr <=  "0000000110000";
		Trees_din <= x"190e000c";
		wait for Clk_period;
		Addr <=  "0000000110001";
		Trees_din <= x"3a0b9804";
		wait for Clk_period;
		Addr <=  "0000000110010";
		Trees_din <= x"ff580115";
		wait for Clk_period;
		Addr <=  "0000000110011";
		Trees_din <= x"c5047c04";
		wait for Clk_period;
		Addr <=  "0000000110100";
		Trees_din <= x"ff6a0115";
		wait for Clk_period;
		Addr <=  "0000000110101";
		Trees_din <= x"00d50115";
		wait for Clk_period;
		Addr <=  "0000000110110";
		Trees_din <= x"00010115";
		wait for Clk_period;
		Addr <=  "0000000110111";
		Trees_din <= x"1a05d508";
		wait for Clk_period;
		Addr <=  "0000000111000";
		Trees_din <= x"d8023604";
		wait for Clk_period;
		Addr <=  "0000000111001";
		Trees_din <= x"003f0115";
		wait for Clk_period;
		Addr <=  "0000000111010";
		Trees_din <= x"ff6f0115";
		wait for Clk_period;
		Addr <=  "0000000111011";
		Trees_din <= x"01720115";
		wait for Clk_period;
		Addr <=  "0000000111100";
		Trees_din <= x"00020208";
		wait for Clk_period;
		Addr <=  "0000000111101";
		Trees_din <= x"01006f04";
		wait for Clk_period;
		Addr <=  "0000000111110";
		Trees_din <= x"00860115";
		wait for Clk_period;
		Addr <=  "0000000111111";
		Trees_din <= x"ff780115";
		wait for Clk_period;
		Addr <=  "0000001000000";
		Trees_din <= x"1603b908";
		wait for Clk_period;
		Addr <=  "0000001000001";
		Trees_din <= x"cd006904";
		wait for Clk_period;
		Addr <=  "0000001000010";
		Trees_din <= x"00840115";
		wait for Clk_period;
		Addr <=  "0000001000011";
		Trees_din <= x"000b0115";
		wait for Clk_period;
		Addr <=  "0000001000100";
		Trees_din <= x"01440115";
		wait for Clk_period;
		Addr <=  "0000001000101";
		Trees_din <= x"1a08a114";
		wait for Clk_period;
		Addr <=  "0000001000110";
		Trees_din <= x"190e000c";
		wait for Clk_period;
		Addr <=  "0000001000111";
		Trees_din <= x"e311c604";
		wait for Clk_period;
		Addr <=  "0000001001000";
		Trees_din <= x"ff5c0169";
		wait for Clk_period;
		Addr <=  "0000001001001";
		Trees_din <= x"26010304";
		wait for Clk_period;
		Addr <=  "0000001001010";
		Trees_din <= x"ff7f0169";
		wait for Clk_period;
		Addr <=  "0000001001011";
		Trees_din <= x"00ae0169";
		wait for Clk_period;
		Addr <=  "0000001001100";
		Trees_din <= x"03052304";
		wait for Clk_period;
		Addr <=  "0000001001101";
		Trees_din <= x"ffa00169";
		wait for Clk_period;
		Addr <=  "0000001001110";
		Trees_din <= x"01230169";
		wait for Clk_period;
		Addr <=  "0000001001111";
		Trees_din <= x"43057708";
		wait for Clk_period;
		Addr <=  "0000001010000";
		Trees_din <= x"4200c304";
		wait for Clk_period;
		Addr <=  "0000001010001";
		Trees_din <= x"00210169";
		wait for Clk_period;
		Addr <=  "0000001010010";
		Trees_din <= x"ff6b0169";
		wait for Clk_period;
		Addr <=  "0000001010011";
		Trees_din <= x"78023e04";
		wait for Clk_period;
		Addr <=  "0000001010100";
		Trees_din <= x"ff9f0169";
		wait for Clk_period;
		Addr <=  "0000001010101";
		Trees_din <= x"d2073a04";
		wait for Clk_period;
		Addr <=  "0000001010110";
		Trees_din <= x"ffa10169";
		wait for Clk_period;
		Addr <=  "0000001010111";
		Trees_din <= x"7c074804";
		wait for Clk_period;
		Addr <=  "0000001011000";
		Trees_din <= x"010f0169";
		wait for Clk_period;
		Addr <=  "0000001011001";
		Trees_din <= x"00490169";
		wait for Clk_period;
		Addr <=  "0000001011010";
		Trees_din <= x"1a08a114";
		wait for Clk_period;
		Addr <=  "0000001011011";
		Trees_din <= x"190e000c";
		wait for Clk_period;
		Addr <=  "0000001011100";
		Trees_din <= x"e311c604";
		wait for Clk_period;
		Addr <=  "0000001011101";
		Trees_din <= x"ff5e01bd";
		wait for Clk_period;
		Addr <=  "0000001011110";
		Trees_din <= x"5e017b04";
		wait for Clk_period;
		Addr <=  "0000001011111";
		Trees_din <= x"ff8601bd";
		wait for Clk_period;
		Addr <=  "0000001100000";
		Trees_din <= x"009901bd";
		wait for Clk_period;
		Addr <=  "0000001100001";
		Trees_din <= x"03052304";
		wait for Clk_period;
		Addr <=  "0000001100010";
		Trees_din <= x"ffa901bd";
		wait for Clk_period;
		Addr <=  "0000001100011";
		Trees_din <= x"00f301bd";
		wait for Clk_period;
		Addr <=  "0000001100100";
		Trees_din <= x"1708c508";
		wait for Clk_period;
		Addr <=  "0000001100101";
		Trees_din <= x"1d004e04";
		wait for Clk_period;
		Addr <=  "0000001100110";
		Trees_din <= x"007301bd";
		wait for Clk_period;
		Addr <=  "0000001100111";
		Trees_din <= x"ff6f01bd";
		wait for Clk_period;
		Addr <=  "0000001101000";
		Trees_din <= x"d2073a04";
		wait for Clk_period;
		Addr <=  "0000001101001";
		Trees_din <= x"ff9e01bd";
		wait for Clk_period;
		Addr <=  "0000001101010";
		Trees_din <= x"f804f804";
		wait for Clk_period;
		Addr <=  "0000001101011";
		Trees_din <= x"00e801bd";
		wait for Clk_period;
		Addr <=  "0000001101100";
		Trees_din <= x"2b089104";
		wait for Clk_period;
		Addr <=  "0000001101101";
		Trees_din <= x"005901bd";
		wait for Clk_period;
		Addr <=  "0000001101110";
		Trees_din <= x"fffd01bd";
		wait for Clk_period;
		Addr <=  "0000001101111";
		Trees_din <= x"1a08a114";
		wait for Clk_period;
		Addr <=  "0000001110000";
		Trees_din <= x"190e000c";
		wait for Clk_period;
		Addr <=  "0000001110001";
		Trees_din <= x"e311c604";
		wait for Clk_period;
		Addr <=  "0000001110010";
		Trees_din <= x"ff600211";
		wait for Clk_period;
		Addr <=  "0000001110011";
		Trees_din <= x"37038404";
		wait for Clk_period;
		Addr <=  "0000001110100";
		Trees_din <= x"ff8e0211";
		wait for Clk_period;
		Addr <=  "0000001110101";
		Trees_din <= x"008b0211";
		wait for Clk_period;
		Addr <=  "0000001110110";
		Trees_din <= x"7d009104";
		wait for Clk_period;
		Addr <=  "0000001110111";
		Trees_din <= x"00af0211";
		wait for Clk_period;
		Addr <=  "0000001111000";
		Trees_din <= x"00050211";
		wait for Clk_period;
		Addr <=  "0000001111001";
		Trees_din <= x"43057708";
		wait for Clk_period;
		Addr <=  "0000001111010";
		Trees_din <= x"5b079f04";
		wait for Clk_period;
		Addr <=  "0000001111011";
		Trees_din <= x"ff780211";
		wait for Clk_period;
		Addr <=  "0000001111100";
		Trees_din <= x"00090211";
		wait for Clk_period;
		Addr <=  "0000001111101";
		Trees_din <= x"b5011004";
		wait for Clk_period;
		Addr <=  "0000001111110";
		Trees_din <= x"ffd30211";
		wait for Clk_period;
		Addr <=  "0000001111111";
		Trees_din <= x"62022a08";
		wait for Clk_period;
		Addr <=  "0000010000000";
		Trees_din <= x"1c00a704";
		wait for Clk_period;
		Addr <=  "0000010000001";
		Trees_din <= x"001d0211";
		wait for Clk_period;
		Addr <=  "0000010000010";
		Trees_din <= x"00d10211";
		wait for Clk_period;
		Addr <=  "0000010000011";
		Trees_din <= x"ffee0211";
		wait for Clk_period;
		Addr <=  "0000010000100";
		Trees_din <= x"1a08a114";
		wait for Clk_period;
		Addr <=  "0000010000101";
		Trees_din <= x"190e000c";
		wait for Clk_period;
		Addr <=  "0000010000110";
		Trees_din <= x"e311c604";
		wait for Clk_period;
		Addr <=  "0000010000111";
		Trees_din <= x"ff62025d";
		wait for Clk_period;
		Addr <=  "0000010001000";
		Trees_din <= x"5b020c04";
		wait for Clk_period;
		Addr <=  "0000010001001";
		Trees_din <= x"ff97025d";
		wait for Clk_period;
		Addr <=  "0000010001010";
		Trees_din <= x"007a025d";
		wait for Clk_period;
		Addr <=  "0000010001011";
		Trees_din <= x"bc03d204";
		wait for Clk_period;
		Addr <=  "0000010001100";
		Trees_din <= x"00a5025d";
		wait for Clk_period;
		Addr <=  "0000010001101";
		Trees_din <= x"0009025d";
		wait for Clk_period;
		Addr <=  "0000010001110";
		Trees_din <= x"1708c508";
		wait for Clk_period;
		Addr <=  "0000010001111";
		Trees_din <= x"ae007204";
		wait for Clk_period;
		Addr <=  "0000010010000";
		Trees_din <= x"004d025d";
		wait for Clk_period;
		Addr <=  "0000010010001";
		Trees_din <= x"ff7b025d";
		wait for Clk_period;
		Addr <=  "0000010010010";
		Trees_din <= x"d2073a04";
		wait for Clk_period;
		Addr <=  "0000010010011";
		Trees_din <= x"ffac025d";
		wait for Clk_period;
		Addr <=  "0000010010100";
		Trees_din <= x"f804f804";
		wait for Clk_period;
		Addr <=  "0000010010101";
		Trees_din <= x"00c0025d";
		wait for Clk_period;
		Addr <=  "0000010010110";
		Trees_din <= x"0029025d";
		wait for Clk_period;
		Addr <=  "0000010010111";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0000010011000";
		Trees_din <= x"1a08a114";
		wait for Clk_period;
		Addr <=  "0000010011001";
		Trees_din <= x"190e000c";
		wait for Clk_period;
		Addr <=  "0000010011010";
		Trees_din <= x"e311c604";
		wait for Clk_period;
		Addr <=  "0000010011011";
		Trees_din <= x"ff6302ad";
		wait for Clk_period;
		Addr <=  "0000010011100";
		Trees_din <= x"2600d004";
		wait for Clk_period;
		Addr <=  "0000010011101";
		Trees_din <= x"ffa102ad";
		wait for Clk_period;
		Addr <=  "0000010011110";
		Trees_din <= x"006602ad";
		wait for Clk_period;
		Addr <=  "0000010011111";
		Trees_din <= x"7902f604";
		wait for Clk_period;
		Addr <=  "0000010100000";
		Trees_din <= x"009402ad";
		wait for Clk_period;
		Addr <=  "0000010100001";
		Trees_din <= x"000802ad";
		wait for Clk_period;
		Addr <=  "0000010100010";
		Trees_din <= x"43057708";
		wait for Clk_period;
		Addr <=  "0000010100011";
		Trees_din <= x"0d008704";
		wait for Clk_period;
		Addr <=  "0000010100100";
		Trees_din <= x"fff302ad";
		wait for Clk_period;
		Addr <=  "0000010100101";
		Trees_din <= x"ff8702ad";
		wait for Clk_period;
		Addr <=  "0000010100110";
		Trees_din <= x"49048b08";
		wait for Clk_period;
		Addr <=  "0000010100111";
		Trees_din <= x"cf03e904";
		wait for Clk_period;
		Addr <=  "0000010101000";
		Trees_din <= x"002d02ad";
		wait for Clk_period;
		Addr <=  "0000010101001";
		Trees_din <= x"00b502ad";
		wait for Clk_period;
		Addr <=  "0000010101010";
		Trees_din <= x"ffe402ad";
		wait for Clk_period;
		Addr <=  "0000010101011";
		Trees_din <= x"170b9914";
		wait for Clk_period;
		Addr <=  "0000010101100";
		Trees_din <= x"1a0acd0c";
		wait for Clk_period;
		Addr <=  "0000010101101";
		Trees_din <= x"3a0b9804";
		wait for Clk_period;
		Addr <=  "0000010101110";
		Trees_din <= x"ff6402f1";
		wait for Clk_period;
		Addr <=  "0000010101111";
		Trees_din <= x"b103a404";
		wait for Clk_period;
		Addr <=  "0000010110000";
		Trees_din <= x"006802f1";
		wait for Clk_period;
		Addr <=  "0000010110001";
		Trees_din <= x"ff9d02f1";
		wait for Clk_period;
		Addr <=  "0000010110010";
		Trees_din <= x"16059504";
		wait for Clk_period;
		Addr <=  "0000010110011";
		Trees_din <= x"ffa302f1";
		wait for Clk_period;
		Addr <=  "0000010110100";
		Trees_din <= x"006a02f1";
		wait for Clk_period;
		Addr <=  "0000010110101";
		Trees_din <= x"e3058d04";
		wait for Clk_period;
		Addr <=  "0000010110110";
		Trees_din <= x"ff9302f1";
		wait for Clk_period;
		Addr <=  "0000010110111";
		Trees_din <= x"78036004";
		wait for Clk_period;
		Addr <=  "0000010111000";
		Trees_din <= x"ffd602f1";
		wait for Clk_period;
		Addr <=  "0000010111001";
		Trees_din <= x"8d04c204";
		wait for Clk_period;
		Addr <=  "0000010111010";
		Trees_din <= x"002202f1";
		wait for Clk_period;
		Addr <=  "0000010111011";
		Trees_din <= x"00b102f1";
		wait for Clk_period;
		Addr <=  "0000010111100";
		Trees_din <= x"170b9914";
		wait for Clk_period;
		Addr <=  "0000010111101";
		Trees_din <= x"1a0acd0c";
		wait for Clk_period;
		Addr <=  "0000010111110";
		Trees_din <= x"3a0b9804";
		wait for Clk_period;
		Addr <=  "0000010111111";
		Trees_din <= x"ff650335";
		wait for Clk_period;
		Addr <=  "0000011000000";
		Trees_din <= x"f802de04";
		wait for Clk_period;
		Addr <=  "0000011000001";
		Trees_din <= x"00540335";
		wait for Clk_period;
		Addr <=  "0000011000010";
		Trees_din <= x"ffa60335";
		wait for Clk_period;
		Addr <=  "0000011000011";
		Trees_din <= x"2a01b104";
		wait for Clk_period;
		Addr <=  "0000011000100";
		Trees_din <= x"00600335";
		wait for Clk_period;
		Addr <=  "0000011000101";
		Trees_din <= x"ffaa0335";
		wait for Clk_period;
		Addr <=  "0000011000110";
		Trees_din <= x"1a039e08";
		wait for Clk_period;
		Addr <=  "0000011000111";
		Trees_din <= x"fe023604";
		wait for Clk_period;
		Addr <=  "0000011001000";
		Trees_din <= x"ff9f0335";
		wait for Clk_period;
		Addr <=  "0000011001001";
		Trees_din <= x"fffb0335";
		wait for Clk_period;
		Addr <=  "0000011001010";
		Trees_din <= x"3a075904";
		wait for Clk_period;
		Addr <=  "0000011001011";
		Trees_din <= x"00080335";
		wait for Clk_period;
		Addr <=  "0000011001100";
		Trees_din <= x"00a50335";
		wait for Clk_period;
		Addr <=  "0000011001101";
		Trees_din <= x"170b9914";
		wait for Clk_period;
		Addr <=  "0000011001110";
		Trees_din <= x"1a096808";
		wait for Clk_period;
		Addr <=  "0000011001111";
		Trees_din <= x"e311c604";
		wait for Clk_period;
		Addr <=  "0000011010000";
		Trees_din <= x"ff660379";
		wait for Clk_period;
		Addr <=  "0000011010001";
		Trees_din <= x"fffe0379";
		wait for Clk_period;
		Addr <=  "0000011010010";
		Trees_din <= x"85081a04";
		wait for Clk_period;
		Addr <=  "0000011010011";
		Trees_din <= x"ff9e0379";
		wait for Clk_period;
		Addr <=  "0000011010100";
		Trees_din <= x"e8039704";
		wait for Clk_period;
		Addr <=  "0000011010101";
		Trees_din <= x"00680379";
		wait for Clk_period;
		Addr <=  "0000011010110";
		Trees_din <= x"00180379";
		wait for Clk_period;
		Addr <=  "0000011010111";
		Trees_din <= x"85058708";
		wait for Clk_period;
		Addr <=  "0000011011000";
		Trees_din <= x"f505c504";
		wait for Clk_period;
		Addr <=  "0000011011001";
		Trees_din <= x"ff9c0379";
		wait for Clk_period;
		Addr <=  "0000011011010";
		Trees_din <= x"00200379";
		wait for Clk_period;
		Addr <=  "0000011011011";
		Trees_din <= x"22034704";
		wait for Clk_period;
		Addr <=  "0000011011100";
		Trees_din <= x"00a20379";
		wait for Clk_period;
		Addr <=  "0000011011101";
		Trees_din <= x"00090379";
		wait for Clk_period;
		Addr <=  "0000011011110";
		Trees_din <= x"3a086610";
		wait for Clk_period;
		Addr <=  "0000011011111";
		Trees_din <= x"850b0108";
		wait for Clk_period;
		Addr <=  "0000011100000";
		Trees_din <= x"ce09c504";
		wait for Clk_period;
		Addr <=  "0000011100001";
		Trees_din <= x"ff6603b5";
		wait for Clk_period;
		Addr <=  "0000011100010";
		Trees_din <= x"ffd403b5";
		wait for Clk_period;
		Addr <=  "0000011100011";
		Trees_din <= x"1a074304";
		wait for Clk_period;
		Addr <=  "0000011100100";
		Trees_din <= x"ffad03b5";
		wait for Clk_period;
		Addr <=  "0000011100101";
		Trees_din <= x"004f03b5";
		wait for Clk_period;
		Addr <=  "0000011100110";
		Trees_din <= x"f8058b0c";
		wait for Clk_period;
		Addr <=  "0000011100111";
		Trees_din <= x"78039704";
		wait for Clk_period;
		Addr <=  "0000011101000";
		Trees_din <= x"fff803b5";
		wait for Clk_period;
		Addr <=  "0000011101001";
		Trees_din <= x"8301fa04";
		wait for Clk_period;
		Addr <=  "0000011101010";
		Trees_din <= x"009d03b5";
		wait for Clk_period;
		Addr <=  "0000011101011";
		Trees_din <= x"003103b5";
		wait for Clk_period;
		Addr <=  "0000011101100";
		Trees_din <= x"ffa203b5";
		wait for Clk_period;
		Addr <=  "0000011101101";
		Trees_din <= x"1a08170c";
		wait for Clk_period;
		Addr <=  "0000011101110";
		Trees_din <= x"3a086604";
		wait for Clk_period;
		Addr <=  "0000011101111";
		Trees_din <= x"ff6703e1";
		wait for Clk_period;
		Addr <=  "0000011110000";
		Trees_din <= x"f8012b04";
		wait for Clk_period;
		Addr <=  "0000011110001";
		Trees_din <= x"005703e1";
		wait for Clk_period;
		Addr <=  "0000011110010";
		Trees_din <= x"ff9403e1";
		wait for Clk_period;
		Addr <=  "0000011110011";
		Trees_din <= x"43057704";
		wait for Clk_period;
		Addr <=  "0000011110100";
		Trees_din <= x"ffb003e1";
		wait for Clk_period;
		Addr <=  "0000011110101";
		Trees_din <= x"8d04c204";
		wait for Clk_period;
		Addr <=  "0000011110110";
		Trees_din <= x"fffc03e1";
		wait for Clk_period;
		Addr <=  "0000011110111";
		Trees_din <= x"009003e1";
		wait for Clk_period;
		Addr <=  "0000011111000";
		Trees_din <= x"3a08660c";
		wait for Clk_period;
		Addr <=  "0000011111001";
		Trees_din <= x"1a08a104";
		wait for Clk_period;
		Addr <=  "0000011111010";
		Trees_din <= x"ff68040d";
		wait for Clk_period;
		Addr <=  "0000011111011";
		Trees_din <= x"01012e04";
		wait for Clk_period;
		Addr <=  "0000011111100";
		Trees_din <= x"0037040d";
		wait for Clk_period;
		Addr <=  "0000011111101";
		Trees_din <= x"ffad040d";
		wait for Clk_period;
		Addr <=  "0000011111110";
		Trees_din <= x"5e036304";
		wait for Clk_period;
		Addr <=  "0000011111111";
		Trees_din <= x"ffb1040d";
		wait for Clk_period;
		Addr <=  "0000100000000";
		Trees_din <= x"dd03ed04";
		wait for Clk_period;
		Addr <=  "0000100000001";
		Trees_din <= x"008e040d";
		wait for Clk_period;
		Addr <=  "0000100000010";
		Trees_din <= x"0007040d";
		wait for Clk_period;
		Addr <=  "0000100000011";
		Trees_din <= x"170b9910";
		wait for Clk_period;
		Addr <=  "0000100000100";
		Trees_din <= x"1a096808";
		wait for Clk_period;
		Addr <=  "0000100000101";
		Trees_din <= x"3f000004";
		wait for Clk_period;
		Addr <=  "0000100000110";
		Trees_din <= x"ffe70439";
		wait for Clk_period;
		Addr <=  "0000100000111";
		Trees_din <= x"ff690439";
		wait for Clk_period;
		Addr <=  "0000100001000";
		Trees_din <= x"db013104";
		wait for Clk_period;
		Addr <=  "0000100001001";
		Trees_din <= x"003e0439";
		wait for Clk_period;
		Addr <=  "0000100001010";
		Trees_din <= x"ffc70439";
		wait for Clk_period;
		Addr <=  "0000100001011";
		Trees_din <= x"85058704";
		wait for Clk_period;
		Addr <=  "0000100001100";
		Trees_din <= x"ffdd0439";
		wait for Clk_period;
		Addr <=  "0000100001101";
		Trees_din <= x"00840439";
		wait for Clk_period;
		Addr <=  "0000100001110";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0000100001111";
		Trees_din <= x"3a086608";
		wait for Clk_period;
		Addr <=  "0000100010000";
		Trees_din <= x"850b0104";
		wait for Clk_period;
		Addr <=  "0000100010001";
		Trees_din <= x"ff6b0461";
		wait for Clk_period;
		Addr <=  "0000100010010";
		Trees_din <= x"00020461";
		wait for Clk_period;
		Addr <=  "0000100010011";
		Trees_din <= x"78039d04";
		wait for Clk_period;
		Addr <=  "0000100010100";
		Trees_din <= x"ffc10461";
		wait for Clk_period;
		Addr <=  "0000100010101";
		Trees_din <= x"8d047c04";
		wait for Clk_period;
		Addr <=  "0000100010110";
		Trees_din <= x"00190461";
		wait for Clk_period;
		Addr <=  "0000100010111";
		Trees_din <= x"00850461";
		wait for Clk_period;
		Addr <=  "0000100011000";
		Trees_din <= x"1a081708";
		wait for Clk_period;
		Addr <=  "0000100011001";
		Trees_din <= x"4308b904";
		wait for Clk_period;
		Addr <=  "0000100011010";
		Trees_din <= x"ff6b047d";
		wait for Clk_period;
		Addr <=  "0000100011011";
		Trees_din <= x"fff0047d";
		wait for Clk_period;
		Addr <=  "0000100011100";
		Trees_din <= x"00034904";
		wait for Clk_period;
		Addr <=  "0000100011101";
		Trees_din <= x"ffd9047d";
		wait for Clk_period;
		Addr <=  "0000100011110";
		Trees_din <= x"007a047d";
		wait for Clk_period;
		Addr <=  "0000100011111";
		Trees_din <= x"3a086608";
		wait for Clk_period;
		Addr <=  "0000100100000";
		Trees_din <= x"67091704";
		wait for Clk_period;
		Addr <=  "0000100100001";
		Trees_din <= x"ff6d04a1";
		wait for Clk_period;
		Addr <=  "0000100100010";
		Trees_din <= x"ffe504a1";
		wait for Clk_period;
		Addr <=  "0000100100011";
		Trees_din <= x"5e036304";
		wait for Clk_period;
		Addr <=  "0000100100100";
		Trees_din <= x"ffc804a1";
		wait for Clk_period;
		Addr <=  "0000100100101";
		Trees_din <= x"7107c804";
		wait for Clk_period;
		Addr <=  "0000100100110";
		Trees_din <= x"001e04a1";
		wait for Clk_period;
		Addr <=  "0000100100111";
		Trees_din <= x"007d04a1";
		wait for Clk_period;
		Addr <=  "0000100101000";
		Trees_din <= x"1709f308";
		wait for Clk_period;
		Addr <=  "0000100101001";
		Trees_din <= x"85088104";
		wait for Clk_period;
		Addr <=  "0000100101010";
		Trees_din <= x"ff6e04bd";
		wait for Clk_period;
		Addr <=  "0000100101011";
		Trees_din <= x"ffe404bd";
		wait for Clk_period;
		Addr <=  "0000100101100";
		Trees_din <= x"8d04ca04";
		wait for Clk_period;
		Addr <=  "0000100101101";
		Trees_din <= x"ffd504bd";
		wait for Clk_period;
		Addr <=  "0000100101110";
		Trees_din <= x"007204bd";
		wait for Clk_period;
		Addr <=  "0000100101111";
		Trees_din <= x"3a086608";
		wait for Clk_period;
		Addr <=  "0000100110000";
		Trees_din <= x"67091704";
		wait for Clk_period;
		Addr <=  "0000100110001";
		Trees_din <= x"ff7104d9";
		wait for Clk_period;
		Addr <=  "0000100110010";
		Trees_din <= x"ffeb04d9";
		wait for Clk_period;
		Addr <=  "0000100110011";
		Trees_din <= x"f802ac04";
		wait for Clk_period;
		Addr <=  "0000100110100";
		Trees_din <= x"006c04d9";
		wait for Clk_period;
		Addr <=  "0000100110101";
		Trees_din <= x"ffdf04d9";
		wait for Clk_period;
		Addr <=  "0000100110110";
		Trees_din <= x"1a081708";
		wait for Clk_period;
		Addr <=  "0000100110111";
		Trees_din <= x"4308b904";
		wait for Clk_period;
		Addr <=  "0000100111000";
		Trees_din <= x"ff7304f5";
		wait for Clk_period;
		Addr <=  "0000100111001";
		Trees_din <= x"fff904f5";
		wait for Clk_period;
		Addr <=  "0000100111010";
		Trees_din <= x"0004f604";
		wait for Clk_period;
		Addr <=  "0000100111011";
		Trees_din <= x"000104f5";
		wait for Clk_period;
		Addr <=  "0000100111100";
		Trees_din <= x"006b04f5";
		wait for Clk_period;
		Addr <=  "0000100111101";
		Trees_din <= x"1a081708";
		wait for Clk_period;
		Addr <=  "0000100111110";
		Trees_din <= x"4308b904";
		wait for Clk_period;
		Addr <=  "0000100111111";
		Trees_din <= x"ff760511";
		wait for Clk_period;
		Addr <=  "0000101000000";
		Trees_din <= x"fffb0511";
		wait for Clk_period;
		Addr <=  "0000101000001";
		Trees_din <= x"0004f604";
		wait for Clk_period;
		Addr <=  "0000101000010";
		Trees_din <= x"00010511";
		wait for Clk_period;
		Addr <=  "0000101000011";
		Trees_din <= x"00650511";
		wait for Clk_period;
		Addr <=  "0000101000100";
		Trees_din <= x"1709f308";
		wait for Clk_period;
		Addr <=  "0000101000101";
		Trees_din <= x"67072f04";
		wait for Clk_period;
		Addr <=  "0000101000110";
		Trees_din <= x"ff7c052d";
		wait for Clk_period;
		Addr <=  "0000101000111";
		Trees_din <= x"ffdf052d";
		wait for Clk_period;
		Addr <=  "0000101001000";
		Trees_din <= x"8d074004";
		wait for Clk_period;
		Addr <=  "0000101001001";
		Trees_din <= x"0001052d";
		wait for Clk_period;
		Addr <=  "0000101001010";
		Trees_din <= x"0061052d";
		wait for Clk_period;
		Addr <=  "0000101001011";
		Trees_din <= x"3a086608";
		wait for Clk_period;
		Addr <=  "0000101001100";
		Trees_din <= x"43057704";
		wait for Clk_period;
		Addr <=  "0000101001101";
		Trees_din <= x"ff7f0549";
		wait for Clk_period;
		Addr <=  "0000101001110";
		Trees_din <= x"ffe10549";
		wait for Clk_period;
		Addr <=  "0000101001111";
		Trees_din <= x"8d065d04";
		wait for Clk_period;
		Addr <=  "0000101010000";
		Trees_din <= x"fffd0549";
		wait for Clk_period;
		Addr <=  "0000101010001";
		Trees_din <= x"005c0549";
		wait for Clk_period;
		Addr <=  "0000101010010";
		Trees_din <= x"1a081708";
		wait for Clk_period;
		Addr <=  "0000101010011";
		Trees_din <= x"71079604";
		wait for Clk_period;
		Addr <=  "0000101010100";
		Trees_din <= x"ff830565";
		wait for Clk_period;
		Addr <=  "0000101010101";
		Trees_din <= x"ffec0565";
		wait for Clk_period;
		Addr <=  "0000101010110";
		Trees_din <= x"5e06eb04";
		wait for Clk_period;
		Addr <=  "0000101010111";
		Trees_din <= x"00130565";
		wait for Clk_period;
		Addr <=  "0000101011000";
		Trees_din <= x"00530565";
		wait for Clk_period;
		Addr <=  "0000101011001";
		Trees_din <= x"3a086604";
		wait for Clk_period;
		Addr <=  "0000101011010";
		Trees_din <= x"ff920579";
		wait for Clk_period;
		Addr <=  "0000101011011";
		Trees_din <= x"cd023404";
		wait for Clk_period;
		Addr <=  "0000101011100";
		Trees_din <= x"004b0579";
		wait for Clk_period;
		Addr <=  "0000101011101";
		Trees_din <= x"00110579";
		wait for Clk_period;
		Addr <=  "0000101011110";
		Trees_din <= x"170b9908";
		wait for Clk_period;
		Addr <=  "0000101011111";
		Trees_din <= x"85063c04";
		wait for Clk_period;
		Addr <=  "0000101100000";
		Trees_din <= x"ff8d058d";
		wait for Clk_period;
		Addr <=  "0000101100001";
		Trees_din <= x"ffec058d";
		wait for Clk_period;
		Addr <=  "0000101100010";
		Trees_din <= x"0048058d";
		wait for Clk_period;
		Addr <=  "0000101100011";
		Trees_din <= x"43057704";
		wait for Clk_period;
		Addr <=  "0000101100100";
		Trees_din <= x"ff9105a1";
		wait for Clk_period;
		Addr <=  "0000101100101";
		Trees_din <= x"78070d04";
		wait for Clk_period;
		Addr <=  "0000101100110";
		Trees_din <= x"fff405a1";
		wait for Clk_period;
		Addr <=  "0000101100111";
		Trees_din <= x"005005a1";
		wait for Clk_period;
		Addr <=  "0000101101000";
		Trees_din <= x"71079604";
		wait for Clk_period;
		Addr <=  "0000101101001";
		Trees_din <= x"ff9f05ad";
		wait for Clk_period;
		Addr <=  "0000101101010";
		Trees_din <= x"003505ad";
		wait for Clk_period;
		Addr <=  "0000101101011";
		Trees_din <= x"43057704";
		wait for Clk_period;
		Addr <=  "0000101101100";
		Trees_din <= x"ff9b05c1";
		wait for Clk_period;
		Addr <=  "0000101101101";
		Trees_din <= x"78070d04";
		wait for Clk_period;
		Addr <=  "0000101101110";
		Trees_din <= x"fff905c1";
		wait for Clk_period;
		Addr <=  "0000101101111";
		Trees_din <= x"004b05c1";
		wait for Clk_period;
		Addr <=  "0000101110000";
		Trees_din <= x"1a081704";
		wait for Clk_period;
		Addr <=  "0000101110001";
		Trees_din <= x"ffac05cd";
		wait for Clk_period;
		Addr <=  "0000101110010";
		Trees_din <= x"003a05cd";
		wait for Clk_period;
		Addr <=  "0000101110011";
		Trees_din <= x"85069204";
		wait for Clk_period;
		Addr <=  "0000101110100";
		Trees_din <= x"ffa905d9";
		wait for Clk_period;
		Addr <=  "0000101110101";
		Trees_din <= x"002e05d9";
		wait for Clk_period;
		Addr <=  "0000101110110";
		Trees_din <= x"3a086604";
		wait for Clk_period;
		Addr <=  "0000101110111";
		Trees_din <= x"ffb205e5";
		wait for Clk_period;
		Addr <=  "0000101111000";
		Trees_din <= x"003305e5";
		wait for Clk_period;
		Addr <=  "0000101111001";
		Trees_din <= x"43057704";
		wait for Clk_period;
		Addr <=  "0000101111010";
		Trees_din <= x"ffae05f1";
		wait for Clk_period;
		Addr <=  "0000101111011";
		Trees_din <= x"002905f1";
		wait for Clk_period;
		Addr <=  "0000101111100";
		Trees_din <= x"71079604";
		wait for Clk_period;
		Addr <=  "0000101111101";
		Trees_din <= x"ffb805fd";
		wait for Clk_period;
		Addr <=  "0000101111110";
		Trees_din <= x"002f05fd";
		wait for Clk_period;
		Addr <=  "0000101111111";
		Trees_din <= x"1a081704";
		wait for Clk_period;
		Addr <=  "0000110000000";
		Trees_din <= x"ffbe0609";
		wait for Clk_period;
		Addr <=  "0000110000001";
		Trees_din <= x"00300609";
		wait for Clk_period;
		Addr <=  "0000110000010";
		Trees_din <= x"78054a04";
		wait for Clk_period;
		Addr <=  "0000110000011";
		Trees_din <= x"ffc10615";
		wait for Clk_period;
		Addr <=  "0000110000100";
		Trees_din <= x"002d0615";
		wait for Clk_period;
		Addr <=  "0000110000101";
		Trees_din <= x"71079604";
		wait for Clk_period;
		Addr <=  "0000110000110";
		Trees_din <= x"ffc30621";
		wait for Clk_period;
		Addr <=  "0000110000111";
		Trees_din <= x"002a0621";
		wait for Clk_period;
		Addr <=  "0000110001000";
		Trees_din <= x"7804aa04";
		wait for Clk_period;
		Addr <=  "0000110001001";
		Trees_din <= x"ffc6062d";
		wait for Clk_period;
		Addr <=  "0000110001010";
		Trees_din <= x"0029062d";
		wait for Clk_period;
		Addr <=  "0000110001011";
		Trees_din <= x"fff60631";
		wait for Clk_period;
		Addr <=  "0000110001100";
		Trees_din <= x"fff60635";
		wait for Clk_period;
		Addr <=  "0000110001101";
		Trees_din <= x"00000007";
		wait for Clk_period;
		Addr <=  "0000110001110";
		Trees_din <= x"fff7063d";
		wait for Clk_period;
		Addr <=  "0000110001111";
		Trees_din <= x"0000001f";
		wait for Clk_period;

        -- Reset valid flag
        Valid_node <= '0';
        wait for Clk_period; 
        
        class_label <= std_logic_vector(to_unsigned(5, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110100010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010011000000";
        wait for Clk_period; 
        Features_din <= "0000010011111100";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000010010001000";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000010101011110";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000010010111100";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010010000000";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010011000010";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000010111101011";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010010001101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010001011101";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010100001111";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001100010111";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001010100110";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000010011110011";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001100001000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010001111011";
        wait for Clk_period; 
        Features_din <= "0000010011010100";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010001100001";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001100101101";
        wait for Clk_period; 
        Features_din <= "0000010011001001";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010010101100";
        wait for Clk_period; 
        Features_din <= "0000010110011111";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000010010011100";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010010100001";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010010111001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001011110111";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010101101001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010010001101";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111010001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010011101110";
        wait for Clk_period; 
        Features_din <= "0000010101010001";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001100101011";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001100011011";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010001110001";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010010100101";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010110011101";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000010010110110";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000010001010000";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010001010101";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010100000111";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010001101111";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001100110010";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001010001000";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000010011000000";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001100100100";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001100101011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010010011001";
        wait for Clk_period; 
        Features_din <= "0000010001110101";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000010011001011";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010100011100";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000010001110100";
        wait for Clk_period; 
        Features_din <= "0000010111001101";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010001111101";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001100101000";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000010010000101";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010101001001";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010010101001";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110001011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001100100110";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010011100001";
        wait for Clk_period; 
        Features_din <= "0000010100111001";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000010001110001";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010001100010";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010001100100";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010110010001";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010011000110";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000001100011010";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001100010111";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010010110000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000000110101011";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000010011111110";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000010010111010";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010010111000";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001100101010";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000010011101000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010011011011";
        wait for Clk_period; 
        Features_din <= "0000010110111010";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000010001100111";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010011111001";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001011111001";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010100010000";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010001101110";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001100110001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110100111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000010010100101";
        wait for Clk_period; 
        Features_din <= "0000010011010011";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000010010101010";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010010000111";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000010010010001";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000010010101110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010010000000";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001100011111";
        wait for Clk_period; 
        Features_din <= "0000010101100000";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010010000010";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001100011100";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010010110110";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010001001101";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "1111111100010110";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000010011001011";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010010000000";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000010010101001";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010010001001";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010011000110";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000010110000110";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010011001110";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010011111101";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010010011011";
        wait for Clk_period; 
        Features_din <= "0000001100110001";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001100101011";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010010010011";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010110001011";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110111110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010011010101";
        wait for Clk_period; 
        Features_din <= "0000010100100111";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010011101101";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000010010001100";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010110001001";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010011000100";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001100100100";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010100100000";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000000110001010";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000010010010110";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010001101110";
        wait for Clk_period; 
        Features_din <= "0000010010001000";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010010110001";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010011110111";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010010010110";
        wait for Clk_period; 
        Features_din <= "0000010110000100";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010010110000";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010011010000";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010100001010";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010001101110";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111010111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010011110110";
        wait for Clk_period; 
        Features_din <= "0000010010100010";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010010001011";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000010010001011";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000010110100001";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010001011011";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010001111101";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010101001000";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "1111111101001001";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000010010111110";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001100111000";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000010010001010";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000010001101111";
        wait for Clk_period; 
        Features_din <= "0000010011110010";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010011100101";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010010001100";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010011001100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000010011010101";
        wait for Clk_period; 
        Features_din <= "0000010110100001";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010001011011";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010011111101";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010011101110";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010101110010";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010010000001";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110001111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010011001011";
        wait for Clk_period; 
        Features_din <= "0000010010111000";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001100010010";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010010000110";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010001111110";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001100100111";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010010101010";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000010001001101";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000010011010010";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001100110010";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000010101010011";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010001111001";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001100101000";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001100100011";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010011100001";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001100101011";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "1111111110011001";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010011100101";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000010010000000";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000010001111101";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001100001011";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001100010111";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000010011010100";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010001011100";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001100100110";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010011000101";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010010110011";
        wait for Clk_period; 
        Features_din <= "0000010110110110";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000010010101001";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010010111011";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010010011110";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001100011110";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010110011101";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000010010110100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001011101111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110110100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010010010010";
        wait for Clk_period; 
        Features_din <= "0000010100000110";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000010010010101";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001100100000";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010010100011";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001100011110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010001101001";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010001100100";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010111100100";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010001100101";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010010101111";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010101001010";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000000101000011";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000010010101101";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010010001000";
        wait for Clk_period; 
        Features_din <= "0000010010100111";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010001100110";
        wait for Clk_period; 
        Features_din <= "0000010001011101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010010001111";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010010000011";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010010011001";
        wait for Clk_period; 
        Features_din <= "0000010101111001";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010011000001";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000010010011001";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010011010100";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010001110101";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010101000010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010001100110";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110111010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010010100001";
        wait for Clk_period; 
        Features_din <= "0000010100100110";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010001110100";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000010011101111";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010011001001";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000010110001101";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001100011100";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010011001111";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000010100000100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000010001100100";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010001110111";
        wait for Clk_period; 
        Features_din <= "0000010010011010";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010010111110";
        wait for Clk_period; 
        Features_din <= "0000010110000110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010010000110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010011000111";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010110010110";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010010010010";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001101111111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010011010010";
        wait for Clk_period; 
        Features_din <= "0000010100101001";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000010010000111";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010010000000";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000010101010111";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000010001111000";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000010011011100";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000000111010100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010011001110";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010010110100";
        wait for Clk_period; 
        Features_din <= "0000010011010110";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010001011101";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010001111000";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010100010100";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000010110001011";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010011010101";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001100010001";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010011001111";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010101110000";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000010001001101";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110011111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001100100111";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010001111000";
        wait for Clk_period; 
        Features_din <= "0000010010110100";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010010000110";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000010010000111";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010001010101";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001100001110";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010001100011";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010010000101";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010010101111";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010101010101";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001100100000";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010011111101";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "1111111011110111";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000010011011101";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000010010100001";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010001011011";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010100000001";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000010101110011";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001100001000";
        wait for Clk_period; 
        Features_din <= "0000010001100011";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010010111000";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010001111101";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001100101000";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010010101111";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010011110110";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110110110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000010011100101";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010010111110";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000010101000111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010010010011";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010011010001";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010001011101";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001100010100";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010011010100";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001100100110";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000000000000101";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000010011100001";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000010001010101";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001100011100";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010001101001";
        wait for Clk_period; 
        Features_din <= "0000010100001111";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000010011001011";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010011101011";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010010101010";
        wait for Clk_period; 
        Features_din <= "0000010110011000";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000010001101111";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001100010111";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010010100100";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001100011011";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010001110010";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000010101010111";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010010010011";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110010100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010011010000";
        wait for Clk_period; 
        Features_din <= "0000010101001010";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000010010010010";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010100011101";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010011000011";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010010011100";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010010111011";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000010111011010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010010110101";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000010001111100";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010001001101";
        wait for Clk_period; 
        Features_din <= "0000000101111000";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000010010110010";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010010000001";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010001001101";
        wait for Clk_period; 
        Features_din <= "0000010010100111";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010011000000";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010011100110";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010001011100";
        wait for Clk_period; 
        Features_din <= "0000010101100101";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001100101011";
        wait for Clk_period; 
        Features_din <= "0000010011100010";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010010001100";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010101011001";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010010001000";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111100101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000010010000011";
        wait for Clk_period; 
        Features_din <= "0000010101100010";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000010010011000";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000010010010100";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010001110000";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010110000001";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010001111110";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001100011100";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000010010111101";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001100010110";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001010000000";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000010011011010";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001100110000";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010010010011";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001011100010";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000010010011011";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000010001011010";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000010011101011";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001100110010";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010011000000";
        wait for Clk_period; 
        Features_din <= "0000010110111011";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000010010010011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010011111100";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010001111100";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001100010101";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010010000111";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010110001100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000010010100111";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111111000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000010100001000";
        wait for Clk_period; 
        Features_din <= "0000010011111111";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000010100000100";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010011010011";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000010001101111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010001110101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010010010110";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010110101000";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010010000110";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001100110001";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010011101111";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000010100000001";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000010010101010";
        wait for Clk_period; 
        Features_din <= "0000010011000110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000010011000100";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000010010000111";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001100110001";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010010000011";
        wait for Clk_period; 
        Features_din <= "0000010101100111";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010001101111";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010001111001";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010010001010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010100110101";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111000101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010010110110";
        wait for Clk_period; 
        Features_din <= "0000010011011111";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000010001100001";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001100101101";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010010000111";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000010011110010";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010001100110";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001100011001";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001100011111";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010010111000";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "1111111010101000";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000010011001001";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001100100000";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001100001111";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000010010101001";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010001101111";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000010010010111";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010001110010";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010011100101";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010010011001";
        wait for Clk_period; 
        Features_din <= "0000010110001001";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001100101000";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001100101001";
        wait for Clk_period; 
        Features_din <= "0000010010000111";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010011001101";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010100100010";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000010001011101";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111100101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010011101011";
        wait for Clk_period; 
        Features_din <= "0000010011011100";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010001100010";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010011010101";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001100101000";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000010001011101";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010010010001";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010110000100";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010010010010";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001100100000";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010011010001";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010011111101";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010010010011";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000010010001100";
        wait for Clk_period; 
        Features_din <= "0000010010001111";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000010010011110";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000010010111001";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000010010010000";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001100101011";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010100001101";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010010100101";
        wait for Clk_period; 
        Features_din <= "0000010111110011";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010001101001";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010010111101";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001100101011";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001100000000";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010010100000";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000010101111010";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000010010100001";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111101010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010011100000";
        wait for Clk_period; 
        Features_din <= "0000010101011000";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010001101001";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000010011011101";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010010110000";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010010001010";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000010111000001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010010100010";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000010001111101";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001100010110";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010011111001";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "1111101101101101";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000010011111000";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000010010010010";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000010010110100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000010010000101";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010010010111";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000010010001110";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010010011000";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010011011010";
        wait for Clk_period; 
        Features_din <= "0000010111100010";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010001101010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010100010101";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001100110000";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010011011000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001100010110";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010100100011";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111000011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010011001110";
        wait for Clk_period; 
        Features_din <= "0000010100110110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010001111100";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000010110110100";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000010001001101";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010001010101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010010001101";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010010010100";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "1111111100010011";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010011011001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001100000110";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001100111000";
        wait for Clk_period; 
        Features_din <= "0000001100101000";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000010011000111";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000010001111100";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010001110101";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001011110010";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000010001100101";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010011000010";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010001011101";
        wait for Clk_period; 
        Features_din <= "0000010111000001";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000010001101001";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010010100110";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010101100100";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110110000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010010010001";
        wait for Clk_period; 
        Features_din <= "0000010101000110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000010011000010";
        wait for Clk_period; 
        Features_din <= "0000001100011101";
        wait for Clk_period; 
        Features_din <= "0000001100100010";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000010001110001";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010001100101";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000010100101111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010010000101";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010100001000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001001011100";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010001101111";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000010010110100";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010001100001";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000010011001111";
        wait for Clk_period; 
        Features_din <= "0000010110111000";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001100100111";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010010010101";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010011000100";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010010001110";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010110101100";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010010111101";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110111010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000010011010011";
        wait for Clk_period; 
        Features_din <= "0000010101110100";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010010110001";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000010010100100";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000001011011100";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010110111011";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000010010000011";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010001010101";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010010001100";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001011111100";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010011100000";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001000101010";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000010011001110";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000010010000011";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010010000010";
        wait for Clk_period; 
        Features_din <= "0000010011011101";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010001011011";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000010011000010";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010011100111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010001110111";
        wait for Clk_period; 
        Features_din <= "0000010101111001";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000010011000110";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010100000101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010010100000";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001100100100";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010101111010";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110111010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010010000000";
        wait for Clk_period; 
        Features_din <= "0000010100011001";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010010111000";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010001111110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010110001010";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010010010011";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010001011010";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010001101010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001100010000";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010001110001";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010100000111";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "1111111011010100";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000010010011110";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001100010110";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010010001011";
        wait for Clk_period; 
        Features_din <= "0000010001110100";
        wait for Clk_period; 
        Features_din <= "0000001100010110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010001101001";
        wait for Clk_period; 
        Features_din <= "0000010010011110";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010010000110";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000010010001011";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000010011100000";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010010101101";
        wait for Clk_period; 
        Features_din <= "0000010101111100";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010010011011";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000010010101000";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000010100001010";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010001111011";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110000100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010010010100";
        wait for Clk_period; 
        Features_din <= "0000010100110001";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010010001111";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010011101101";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000010010001110";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001100011110";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010011011000";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001100010110";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010101101110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010001100010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001100110000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010001100011";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001100111000";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010011011111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000000100101010";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010010111000";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010001011011";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010010001000";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001100110001";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010100101111";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000010001111101";
        wait for Clk_period; 
        Features_din <= "0000010110101010";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010010000011";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010011000100";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010010110101";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010100111100";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010010111110";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110110010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010010100101";
        wait for Clk_period; 
        Features_din <= "0000010011010111";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010001100100";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000010010110100";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000010001111001";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010001100011";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000010110011110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010010001000";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010010001011";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010010000000";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001100101001";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000010011111001";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000000001010000";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000010010100010";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010001110111";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000010010001000";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010011000111";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000010110101011";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000010010000000";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010010101111";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000010010100011";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010110010010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000010011001101";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110101111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010011010011";
        wait for Clk_period; 
        Features_din <= "0000010100100111";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010010110000";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010001110010";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010010000010";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010010000111";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000010110110000";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010010001000";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010010000100";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001011111101";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000010011010110";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000010010011100";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000010010011111";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010010001011";
        wait for Clk_period; 
        Features_din <= "0000010001100111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001100101010";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000010011001101";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000010001110100";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010011010010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010001111000";
        wait for Clk_period; 
        Features_din <= "0000010111100111";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000010010010011";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010001111000";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001011011100";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001100100100";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010011110110";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110111101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010010000010";
        wait for Clk_period; 
        Features_din <= "0000010100011000";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010010000000";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010010110011";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010010010001";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010001110000";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001100111000";
        wait for Clk_period; 
        Features_din <= "0000010110011101";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010001111011";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010010000110";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010001110000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001011111000";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001100101000";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001100011111";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010010110101";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001100010111";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010011011111";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001100000010";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010010100001";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010001111101";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010011111110";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010011000001";
        wait for Clk_period; 
        Features_din <= "0000010110110100";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000010010100101";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000010010010010";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010010010101";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001100011001";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010110100111";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010010011001";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111100100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000010010100110";
        wait for Clk_period; 
        Features_din <= "0000010011111011";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010010001001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000010010111011";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000010010001100";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001100101000";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010010110001";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010110111101";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010001011011";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010010100110";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001100100100";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010011110010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000000011110010";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000010100000010";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000010010011000";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000010001111001";
        wait for Clk_period; 
        Features_din <= "0000010010101011";
        wait for Clk_period; 
        Features_din <= "0000001100100111";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010010010110";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010010000000";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010010101011";
        wait for Clk_period; 
        Features_din <= "0000010111010001";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001100011101";
        wait for Clk_period; 
        Features_din <= "0000010001110100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010011001000";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010001011011";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001100100000";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010010000010";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010100110011";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(3, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111111001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010011101001";
        wait for Clk_period; 
        Features_din <= "0000010100100000";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010001100001";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010010111001";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000010010010010";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000010010110011";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000010110000010";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010010001110";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010010000000";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010011101111";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000000001011100";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010010100010";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010010001100";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010010000100";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010010000000";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010011000111";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010010010100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000010110111001";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010010011101";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001100010101";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010011000100";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001100111000";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010100110101";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010010100100";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110000001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010100100000";
        wait for Clk_period; 
        Features_din <= "0000010011110010";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010010011001";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000010100000100";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000010010001111";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001100000111";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010001011011";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010010101011";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010001110101";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001100100000";
        wait for Clk_period; 
        Features_din <= "0000010101100101";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001100000001";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010001010101";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010010010101";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000010010001010";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000010001110111";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010010010000";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001100011010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010011110010";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010010110001";
        wait for Clk_period; 
        Features_din <= "0000010110111011";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000010010001111";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010010011000";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010010011011";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001100011100";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010110000001";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010010100101";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001100010001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110011100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010010100010";
        wait for Clk_period; 
        Features_din <= "0000010101100111";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010001110101";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000010100001111";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010010101000";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010010100011";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000010110110101";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010010010001";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010001110000";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000010100111111";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000010011001101";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010010010011";
        wait for Clk_period; 
        Features_din <= "0000010011010010";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000010001110010";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000010010010010";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010011001000";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010010111000";
        wait for Clk_period; 
        Features_din <= "0000010110011010";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000010001111011";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010011010101";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010010100010";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001100110001";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010001100011";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000010100010101";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010010010101";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111001100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010010100010";
        wait for Clk_period; 
        Features_din <= "0000010011100111";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010001111110";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000010010100010";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010010011011";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000010110100111";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000010010001110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010001100010";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010001100011";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001100110010";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010101011011";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001000110101";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000010011101010";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001100001111";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000010010110101";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010001010000";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010001110010";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000010011001101";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010010000011";
        wait for Clk_period; 
        Features_din <= "0000010110000001";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010001101110";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010010010000";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001100100110";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010101000001";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010001101001";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110010101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010100010111";
        wait for Clk_period; 
        Features_din <= "0000010101100101";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010001100110";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010011010001";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010010001100";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001011111111";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000010001111100";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010010110001";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000010110001010";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010001010101";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010010100110";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "1111111101110111";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010001001101";
        wait for Clk_period; 
        Features_din <= "0000010011010011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010001101001";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000010010100011";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001100111000";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010001010101";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001100100010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010011001000";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001100001111";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010001111101";
        wait for Clk_period; 
        Features_din <= "0000010111011111";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001100101000";
        wait for Clk_period; 
        Features_din <= "0000010010111001";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000010010100100";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010010011110";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010110010001";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010010110001";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111010110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000010110100101";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001100100110";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010100011000";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000010010010110";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010011010101";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010001011010";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000010111001101";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010001110111";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010001110101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010001111101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "1111111001100010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000010011001111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010010001001";
        wait for Clk_period; 
        Features_din <= "0000010011001110";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010010010110";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010010011010";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010010101100";
        wait for Clk_period; 
        Features_din <= "0000010101110101";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000010010000010";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010010101010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010010010000";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010010110000";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010100110010";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010001100100";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001100010011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110100111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010010100010";
        wait for Clk_period; 
        Features_din <= "0000010011111001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010010011010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010010101101";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000010100110101";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000010010011010";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010010011000";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000010011000111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "1111111000001110";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010010110001";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000010010110001";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010010001001";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010010010001";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000010010000010";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001100001111";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010010100001";
        wait for Clk_period; 
        Features_din <= "0000010110100011";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001100011001";
        wait for Clk_period; 
        Features_din <= "0000010010001111";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000010010111011";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001100101011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010010110000";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010010100001";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000010110100000";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010010100010";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110110111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010011000011";
        wait for Clk_period; 
        Features_din <= "0000010011010101";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010011000111";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000010010001000";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010001100001";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000010010100010";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010100011101";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010010001100";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010010101011";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010010001011";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010011000100";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001100100000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001001101111";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000010010110001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000010001100110";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010100110101";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001100101001";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000010010110110";
        wait for Clk_period; 
        Features_din <= "0000010111111001";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010100011001";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010010111011";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001011111111";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010001010101";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010101010011";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010001001101";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001101101011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000010011010101";
        wait for Clk_period; 
        Features_din <= "0000010011001000";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010010011011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010010001101";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001100001111";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000010010100001";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000010101011010";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001100101101";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010001001101";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001011111111";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010011100010";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "1111111110101111";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000010011011111";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001011110010";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010010001100";
        wait for Clk_period; 
        Features_din <= "0000010010001000";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010001100001";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000010010111111";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010011001010";
        wait for Clk_period; 
        Features_din <= "0000010110100011";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        Features_din <= "0000010010100001";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001100110010";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010001111001";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010010001100";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010110001110";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010010001100";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111010111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010100001110";
        wait for Clk_period; 
        Features_din <= "0000010011000111";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010001011010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000010011011110";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010010100011";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001100010110";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000010001110001";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010011000000";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010010011110";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000010100100011";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010001111001";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000001100001010";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000000100001110";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010011010101";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010001110000";
        wait for Clk_period; 
        Features_din <= "0000010011111011";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000010001111101";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001100110010";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001100011101";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010010001110";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000010101011110";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000010010101010";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010010001010";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010011000010";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010010010100";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010101011101";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110110010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000010010111010";
        wait for Clk_period; 
        Features_din <= "0000010100111101";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000010011000000";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010011000101";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001011110100";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010001111100";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010010000111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010100100000";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010010010110";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010001101110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001100101101";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001100111000";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010001001101";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010011001100";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001010110000";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000010011101011";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001100100100";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010001100100";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010010111110";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000010110011100";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010010110100";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010010011011";
        wait for Clk_period; 
        Features_din <= "0000001100100000";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010101011100";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010010101000";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110111101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010010000110";
        wait for Clk_period; 
        Features_din <= "0000010101100010";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010010000010";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010010010110";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010010000000";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010011010011";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001100000000";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000010001110101";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010010110011";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001100011101";
        wait for Clk_period; 
        Features_din <= "0000010110001100";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010001111001";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010011001111";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010001001101";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000000111100011";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000010011100011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001010111110";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010001011011";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000010010101100";
        wait for Clk_period; 
        Features_din <= "0000010110011101";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010011111111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001100110000";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010010111010";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010101101100";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010010100001";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111100011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010010110100";
        wait for Clk_period; 
        Features_din <= "0000010100010111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010001010101";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000010010100000";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010101101010";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000010001100001";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010010111110";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001001101000";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000010001110000";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010001011101";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010010000010";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000010001010000";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001100111000";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000010010011110";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000010010110010";
        wait for Clk_period; 
        Features_din <= "0000010110011000";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001100101010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010001110111";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010001111100";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010100100100";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010010011100";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111001110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010011000010";
        wait for Clk_period; 
        Features_din <= "0000010011101111";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010010011100";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001100010000";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010010100001";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000010111001101";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010010000110";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010001100101";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000000101001001";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000010010101001";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010001111000";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001100110010";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000010001110000";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000010001111001";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010011011010";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010010010011";
        wait for Clk_period; 
        Features_din <= "0000010110101010";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010001111000";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001100011111";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010010000011";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010010000010";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010110001111";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000010010001101";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110111001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010100011001";
        wait for Clk_period; 
        Features_din <= "0000010100100100";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000010011110001";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001100100000";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000010010001110";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000010001101111";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010010011000";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010101111110";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010001111011";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010001010000";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001100001001";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010101001000";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010001011100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000000000010001";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000010010001000";
        wait for Clk_period; 
        Features_din <= "0000010011100101";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010001010101";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001011111111";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000010100000000";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000010010100111";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010010111010";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010010001110";
        wait for Clk_period; 
        Features_din <= "0000010101110001";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000010001011101";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001100110010";
        wait for Clk_period; 
        Features_din <= "0000010010110011";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010011011101";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010011010010";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010010100111";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010110100011";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010001110010";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111000010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000010011001011";
        wait for Clk_period; 
        Features_din <= "0000010100100000";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010011000101";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010010100000";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010010001111";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010010011011";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000010110000001";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001100100100";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010100100001";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "1111110111100000";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000010011010101";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000010010001010";
        wait for Clk_period; 
        Features_din <= "0000010010010000";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010010001011";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010100000101";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010010101011";
        wait for Clk_period; 
        Features_din <= "0000010110100000";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000010010011111";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010001101010";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010001101001";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010100110110";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001100011011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110100011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010010100000";
        wait for Clk_period; 
        Features_din <= "0000010101010110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000010010000110";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000010010011001";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010010111001";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010010000110";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000010011011001";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010111010100";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010001011010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010001011101";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010100000110";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001000110100";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000010100000001";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001100100110";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000010010001101";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000010011100100";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010001100010";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010100101101";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000010011000010";
        wait for Clk_period; 
        Features_din <= "0000010111000111";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010010100001";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001100010000";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000010011000101";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010101001001";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010010000101";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001101110011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010010110101";
        wait for Clk_period; 
        Features_din <= "0000010101101000";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010001101110";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010001011011";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010010010001";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010110011010";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000010011000001";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001100101010";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000010010001001";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000010010110100";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000010010100101";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010001100001";
        wait for Clk_period; 
        Features_din <= "0000010011100111";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010011100100";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001100000111";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010011000001";
        wait for Clk_period; 
        Features_din <= "0000010110101010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010010001001";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010100011111";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010010011111";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010100111110";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010001011100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111010000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000010010010101";
        wait for Clk_period; 
        Features_din <= "0000010110000001";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000010100110011";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010001110010";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000010111001110";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010001010101";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000010011000000";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010010011001";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010011000111";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "1111111010000010";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010001111000";
        wait for Clk_period; 
        Features_din <= "0000010011000110";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010010101111";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010010101000";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010010100110";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010010011110";
        wait for Clk_period; 
        Features_din <= "0000010111000110";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010100010111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001100010100";
        wait for Clk_period; 
        Features_din <= "0000001100001110";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000010001101111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010101111101";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000010010101001";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111101001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010011111111";
        wait for Clk_period; 
        Features_din <= "0000010100010011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010001011100";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001100010001";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010010010000";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001100110010";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010001100110";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001011101010";
        wait for Clk_period; 
        Features_din <= "0000010101110110";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010011010111";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010010010001";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001100000001";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001100011100";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010011100011";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001010000101";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000010010110001";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000010011010001";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010010011011";
        wait for Clk_period; 
        Features_din <= "0000010001101010";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000010010101000";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010100010100";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010011010101";
        wait for Clk_period; 
        Features_din <= "0000010101010001";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000010011011011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000010011000001";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001011101010";
        wait for Clk_period; 
        Features_din <= "0000001011110100";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010001110111";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000010101010011";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010010000010";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111001101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010011111001";
        wait for Clk_period; 
        Features_din <= "0000010101001010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001100110001";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010100001100";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000010001100010";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001100101101";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010010001000";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010111000000";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010011000110";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010010011011";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001100011110";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010011100000";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001010110100";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000010001100111";
        wait for Clk_period; 
        Features_din <= "0000010011111101";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010010010111";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000010010011010";
        wait for Clk_period; 
        Features_din <= "0000010010001111";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010001110010";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000010011001111";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010001101110";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010001101110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010010100001";
        wait for Clk_period; 
        Features_din <= "0000010110100000";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010100011001";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001100000111";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010001100010";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001100100011";
        wait for Clk_period; 
        Features_din <= "0000001100000101";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010110000000";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110111100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010100010001";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010001101001";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010010000011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000010100101101";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000010010000110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010010001010";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010001011101";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000010110000010";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010010000100";
        wait for Clk_period; 
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010011110101";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001001011000";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000010010010000";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000010001100010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001100101010";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000010001101001";
        wait for Clk_period; 
        Features_din <= "0000001100101001";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000010010010001";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001100100000";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010011100101";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000001100101010";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010011010010";
        wait for Clk_period; 
        Features_din <= "0000010110110000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001011111011";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010001111101";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010011001111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001011111111";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010101100100";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000010011010011";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001100110000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110110011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010011001011";
        wait for Clk_period; 
        Features_din <= "0000010100011100";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000010001110100";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010001100011";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000010011010100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001100001010";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000010101011101";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010010010101";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001100100110";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000010010010001";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001100100110";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000010011100100";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000010001110101";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010010101001";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010011110111";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010010100111";
        wait for Clk_period; 
        Features_din <= "0000010110100010";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010010011001";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010011010011";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010001110010";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000010001011010";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010101111011";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010010001101";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001101111001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010010101010";
        wait for Clk_period; 
        Features_din <= "0000010100011111";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000010011100111";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010010111010";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000010110010000";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010010101010";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010001011101";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001100100011";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010001100110";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010011111001";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001100001000";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000010011101000";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000010011000010";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010001011100";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010011000011";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000010010111110";
        wait for Clk_period; 
        Features_din <= "0000010110010111";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010100000101";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010010001001";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010110001000";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110101000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010010101111";
        wait for Clk_period; 
        Features_din <= "0000010011010110";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001100100010";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000010011010010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010001111001";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010011000110";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010001010101";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010101001011";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010010010011";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010001111110";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001100100111";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000010001010101";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001001001101";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010011111001";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001100100100";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010001110101";
        wait for Clk_period; 
        Features_din <= "0000010010100011";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010010000101";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010010101011";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000010110010111";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010001110100";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000010101010110";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110100101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010100000111";
        wait for Clk_period; 
        Features_din <= "0000010110100100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010001100101";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010011010100";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010011100000";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001100110010";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010010001110";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010001100111";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010010011011";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010101010100";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001100100100";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010001100101";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010011111100";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000010011101001";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000010010000001";
        wait for Clk_period; 
        Features_din <= "0000010100010000";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010010011001";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010010101010";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010010001001";
        wait for Clk_period; 
        Features_din <= "0000010101010110";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000010011001101";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000010011110011";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010011001100";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010101101001";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010010110110";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110101011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000010011010011";
        wait for Clk_period; 
        Features_din <= "0000010011110100";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010011100000";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000010010101000";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000010001010000";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000010011111111";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001100100000";
        wait for Clk_period; 
        Features_din <= "0000010101010110";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010010001111";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000010001100011";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010011000111";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001100010011";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "1111101111001111";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000010011101101";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000010010110001";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010010001111";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001100011010";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000010010100100";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000010010010100";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000010011100100";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010010000010";
        wait for Clk_period; 
        Features_din <= "0000010110000000";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000010010001101";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001100100010";
        wait for Clk_period; 
        Features_din <= "0000001100001010";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010010010110";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010101110100";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010010000100";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110101010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010011001111";
        wait for Clk_period; 
        Features_din <= "0000010100111010";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000010001101010";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000010011001011";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000010010111100";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000010010011111";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000010101100111";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010010001011";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010001100011";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001100100000";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000010011011000";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010001010101";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000000100011011";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000010100001110";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010010100011";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010001100011";
        wait for Clk_period; 
        Features_din <= "0000010001010101";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010010101101";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001100011110";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010001111100";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010010100001";
        wait for Clk_period; 
        Features_din <= "0000010101001011";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010010001101";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010010100110";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001100011110";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010101101111";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010010001001";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110101101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010011010001";
        wait for Clk_period; 
        Features_din <= "0000010100000000";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001100010010";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000010011100000";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000010010001110";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001100000000";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010010010111";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "0000010110010110";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000010001100011";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010010110101";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000000110101001";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000010010111100";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010001110101";
        wait for Clk_period; 
        Features_din <= "0000010010100010";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000010010101100";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001100011100";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010001111101";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001100010010";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010011100100";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010010101000";
        wait for Clk_period; 
        Features_din <= "0000010111101100";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010010111011";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001100010100";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001100100100";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010010110001";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001100010010";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010101100000";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010010101111";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110000001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010010001010";
        wait for Clk_period; 
        Features_din <= "0000010100111001";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000010010000100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001100010100";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010010010010";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000010110110111";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010001101111";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010010010010";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000010010001010";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001100011001";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001100101000";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001100101101";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001100000100";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001011111001";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000010011101111";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001100011011";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000010010001110";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010001100110";
        wait for Clk_period; 
        Features_din <= "0000010010000010";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001100011111";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000010010010101";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000010011110101";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001011010101";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010010000101";
        wait for Clk_period; 
        Features_din <= "0000010111011100";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010010101100";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010010001000";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000001100011001";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010101010000";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001100101011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110111000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010010111111";
        wait for Clk_period; 
        Features_din <= "0000010100110011";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000010011011001";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010001110101";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000010001101010";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010110010001";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000010010000111";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000010010110011";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010010101000";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010100111011";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000000111111111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000010011100110";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000010001111001";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010001011100";
        wait for Clk_period; 
        Features_din <= "0000010011100100";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010010000000";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010001111100";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000010010110110";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000010010000000";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010010010011";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000010001111101";
        wait for Clk_period; 
        Features_din <= "0000010110000000";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010011001100";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010011001011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010010100010";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010101001010";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010001111100";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(2, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000010000000110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010100000011";
        wait for Clk_period; 
        Features_din <= "0000010011111111";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000010001100101";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010100010010";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010001100100";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010101110000";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010010011111";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001100001011";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010001110101";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010100011000";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000010001100011";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000010010000101";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010010000011";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010011000010";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000010001110010";
        wait for Clk_period; 
        Features_din <= "0000010001110000";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010010101000";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000010111011100";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010010011110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010011011100";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010011011111";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010010111111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(3, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110110101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000010010000011";
        wait for Clk_period; 
        Features_din <= "0000010101001111";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010010000100";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010001011101";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000010011001001";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010010000001";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000010001100110";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010001100001";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010010010001";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010101000111";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001100101000";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000010100000011";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001001111001";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010010011010";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010010011001";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001100110000";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010001011100";
        wait for Clk_period; 
        Features_din <= "0000010011100001";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000010001111011";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010010011111";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010100010010";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000010111011000";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010010011001";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001011111101";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010010101111";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010101111111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010010110001";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110010010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000010100000001";
        wait for Clk_period; 
        Features_din <= "0000010011001011";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010001110000";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000010010011010";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000010011001110";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001100101101";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001100011111";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010011010101";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010101011110";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001011111111";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001100101001";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000010010001010";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010001101111";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010011011100";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001001110011";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000010010100010";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010001010101";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010010010000";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010010001100";
        wait for Clk_period; 
        Features_din <= "0000010010000010";
        wait for Clk_period; 
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010011001010";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010011011111";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010010011000";
        wait for Clk_period; 
        Features_din <= "0000010110000000";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001100100010";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000010010100100";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010010100001";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001100101001";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001100101011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010010000111";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001100100011";
        wait for Clk_period; 
        Features_din <= "0000001100010111";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000010010100110";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010100111101";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000010010111010";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111001100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000010011101010";
        wait for Clk_period; 
        Features_din <= "0000010011011011";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000010010100101";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000010010010010";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000001100110001";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010001110010";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010011011111";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010101111011";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010010000111";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010011001010";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010001011010";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "1111111101100101";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010011000010";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000010001111110";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000010010000001";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010011000011";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000010010100111";
        wait for Clk_period; 
        Features_din <= "0000010110011001";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010001101111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010010111111";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010011000000";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000010110000001";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000010010101001";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110010111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010011000100";
        wait for Clk_period; 
        Features_din <= "0000010101101001";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000010010000110";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000010001111101";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010010010010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010111000001";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001100110001";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010010000011";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001100101000";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010011111011";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000010011101011";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010001100011";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001011111111";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000010011110100";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010010100001";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010010010001";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010010101011";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010011101010";
        wait for Clk_period; 
        Features_din <= "0000010111001000";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010001100010";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010100000100";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010010100011";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001100011101";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010100001111";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010010001111";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(3, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110000010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "0000010100001110";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000010001111101";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010001011100";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000010011010100";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010010100111";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010001110000";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010001111001";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010100101110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000010010000110";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010100110111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "1111110101101100";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001100101010";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010001011010";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010010110010";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010011000010";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000010110010100";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010010111110";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010011001010";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010011101001";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010001010000";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010101101111";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110001110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010010111100";
        wait for Clk_period; 
        Features_din <= "0000010100110011";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010001010101";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010001110001";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000010011101011";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010001011100";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010010101011";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001100101010";
        wait for Clk_period; 
        Features_din <= "0000010110000000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010010101011";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010001011011";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010001100111";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010010101011";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001000011010";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000010011111101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000010010000011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001100100011";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010010001111";
        wait for Clk_period; 
        Features_din <= "0000010010101000";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010001100001";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000010010111101";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001100101011";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000010010101011";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010010101001";
        wait for Clk_period; 
        Features_din <= "0000010111110001";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000010011010001";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010100110111";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010010000100";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010110011010";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010001010000";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110010111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000010011010011";
        wait for Clk_period; 
        Features_din <= "0000010101100100";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010001100100";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010010000001";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000010011111010";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010001110001";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001100110000";
        wait for Clk_period; 
        Features_din <= "0000010110101011";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000010011000100";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010001011010";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010011100100";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001010100111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010011101000";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000010010000111";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010001111110";
        wait for Clk_period; 
        Features_din <= "0000010010000101";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010010000011";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010010101111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010010000010";
        wait for Clk_period; 
        Features_din <= "0000010110010111";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010010111000";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010010111100";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001100011010";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010101101110";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010011000111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001101100110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010011011001";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010010101111";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010010010111";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001100011101";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010011001111";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000010010010000";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010100110110";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010010011010";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000010001100101";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001100000110";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010001111000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000000101110011";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010011010100";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001100011100";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000010010101010";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000010010000010";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001100110000";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010100000101";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000010001100100";
        wait for Clk_period; 
        Features_din <= "0000011000000000";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010011010011";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010010010100";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000010001001101";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010101011110";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110101110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010010010001";
        wait for Clk_period; 
        Features_din <= "0000010101101001";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010001100111";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000010100001110";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000010010000111";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010010010101";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000010110010001";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010001011101";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001100001000";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010001011011";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010100110111";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000010011110010";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010001100001";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010001011011";
        wait for Clk_period; 
        Features_din <= "0000010010100101";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000010010100000";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010010100101";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010011000011";
        wait for Clk_period; 
        Features_din <= "0000010110100100";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010100010000";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010010001100";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000001100010001";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010001110010";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000010101101101";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010010011101";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001100101101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111101111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010010111101";
        wait for Clk_period; 
        Features_din <= "0000010011010111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000010001110000";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001100011100";
        wait for Clk_period; 
        Features_din <= "0000010101011000";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010010010110";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010010101011";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010001111000";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001100001001";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010011110110";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "1111110100110010";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010001010101";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010010001011";
        wait for Clk_period; 
        Features_din <= "0000010001111011";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000010010001111";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010011110110";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010010101100";
        wait for Clk_period; 
        Features_din <= "0000010110010111";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001100100100";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001100101101";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001100010100";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000010010011100";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001100011011";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001100100111";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001011010001";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010010011011";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010100111001";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010010010111";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111010001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000010100001110";
        wait for Clk_period; 
        Features_din <= "0000010011011000";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010001100101";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010011111110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000010010010110";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001100010101";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010010001000";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010010011001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000010101111111";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010001111001";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001100011110";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010011110111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000000110011000";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000010011110000";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010001001101";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010010001000";
        wait for Clk_period; 
        Features_din <= "0000010010100000";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000010001111011";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010010011111";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001100101001";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000010010101001";
        wait for Clk_period; 
        Features_din <= "0000010101110010";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010010100110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010010000011";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001100100011";
        wait for Clk_period; 
        Features_din <= "0000001100101101";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010101111111";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110101110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010011010001";
        wait for Clk_period; 
        Features_din <= "0000010011010001";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010010100001";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010001101110";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010010011111";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000010101000100";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000001100001111";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010001110000";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010100011000";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000000100110001";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000010011011010";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010001110000";
        wait for Clk_period; 
        Features_din <= "0000010010001111";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010010001110";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010010101000";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010001100100";
        wait for Clk_period; 
        Features_din <= "0000010110100110";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001100001000";
        wait for Clk_period; 
        Features_din <= "0000010001110001";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010010001010";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010001100001";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010001100100";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000010110010011";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010010011001";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001100011110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110010101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010011110111";
        wait for Clk_period; 
        Features_din <= "0000010100101101";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010010000101";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000010011010000";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000010001110111";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000010110101000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000010010001000";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000010010101000";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001100101011";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001100100100";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010010100110";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000000110011110";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000010100000100";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001100011001";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010001010000";
        wait for Clk_period; 
        Features_din <= "0000010011010101";
        wait for Clk_period; 
        Features_din <= "0000001100110010";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010011111110";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010011000111";
        wait for Clk_period; 
        Features_din <= "0000010101001000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001100110010";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010001100001";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010011000010";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010010000101";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000010010010101";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010101100100";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001100100110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110101000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010011101010";
        wait for Clk_period; 
        Features_din <= "0000010100110111";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000010011001101";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010010100111";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000010001100001";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010001110001";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000010110011111";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001100110000";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001100011001";
        wait for Clk_period; 
        Features_din <= "0000001100011110";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000010100000010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "1111111011111000";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000010011101111";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010010000101";
        wait for Clk_period; 
        Features_din <= "0000010010110011";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010001010000";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000010010010011";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001100000011";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010011100111";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001100110000";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010001111001";
        wait for Clk_period; 
        Features_din <= "0000010101011011";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001100100111";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001100001100";
        wait for Clk_period; 
        Features_din <= "0000010010101011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010011001111";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000010010011100";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010001111000";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010101011001";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010010011110";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111100100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "0000010100111111";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010010000001";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010001010101";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000010100000011";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000010010110101";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010001110001";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010010000111";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000010110110101";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000010001111100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010001011100";
        wait for Clk_period; 
        Features_din <= "0000001100001110";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001100110001";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010100100011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010001101111";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010010111011";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000010011000000";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010001100110";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001100100100";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000010010000000";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001100000011";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010001011101";
        wait for Clk_period; 
        Features_din <= "0000010011101111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010010001100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010001110111";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000010010011100";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010011110110";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010001110010";
        wait for Clk_period; 
        Features_din <= "0000010110011101";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010011100111";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010010111101";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001100110000";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010001110100";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010100111010";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010010100000";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110010011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010010101110";
        wait for Clk_period; 
        Features_din <= "0000010100011100";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001011101111";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001100111000";
        wait for Clk_period; 
        Features_din <= "0000001100110000";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001100101000";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010011001111";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010101011110";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010010101011";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000010010010000";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001100101101";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001100010001";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000010010011011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000010011111100";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000010010110101";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010010100111";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010010110100";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001100000101";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010010110011";
        wait for Clk_period; 
        Features_din <= "0000010110010111";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000010001100010";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010010110000";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000010101011111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010010011100";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001100001011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001101110101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010100001001";
        wait for Clk_period; 
        Features_din <= "0000010100111011";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010010101010";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000010011010001";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010010100010";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000010010001001";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010101100101";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010010101010";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010010101101";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010001110111";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001011111111";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010011101111";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001100010101";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000010010000100";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000010011110100";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000010001100001";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010011000110";
        wait for Clk_period; 
        Features_din <= "0000010011010011";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010001110101";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010010011000";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010010110101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000010101010011";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000010010101001";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010010110001";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001100101011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010010100101";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010101101110";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010001011101";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110100000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010011010011";
        wait for Clk_period; 
        Features_din <= "0000010100101111";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000010010101011";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000010011010010";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000010010010101";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010010111011";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010001100110";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010011111111";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010001110000";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010001111100";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010011000101";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001100101101";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010001011100";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010010100111";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010010001010";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010010111000";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010010001110";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001100100110";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000010010000101";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010011000001";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000010011011100";
        wait for Clk_period; 
        Features_din <= "0000010110111000";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010010100100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010011011111";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010010001110";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001100111000";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010010110000";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010110001000";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010010100110";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111001000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010100001010";
        wait for Clk_period; 
        Features_din <= "0000010100000101";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010001110010";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010100101111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010010111101";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010111011011";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000010001110100";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000010001011100";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001100011011";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001100001110";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000010010010000";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001010000111";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010010010111";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000010001110100";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000010010101000";
        wait for Clk_period; 
        Features_din <= "0000010010110011";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010001100001";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010010100111";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001100100010";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010011011111";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000010001101010";
        wait for Clk_period; 
        Features_din <= "0000010111000000";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010010001100";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010010101001";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001100110010";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010001111000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010101001101";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111111001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010001101111";
        wait for Clk_period; 
        Features_din <= "0000010101100100";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010001001101";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010001010000";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010010100000";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001100110000";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010001111100";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010111010000";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010001110001";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001100000111";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010010100000";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001000000010";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000010100010010";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000010001110000";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010010011110";
        wait for Clk_period; 
        Features_din <= "0000010010100100";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010001110111";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010010010111";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010010111110";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010010011101";
        wait for Clk_period; 
        Features_din <= "0000010101011110";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010011001010";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010011010011";
        wait for Clk_period; 
        Features_din <= "0000001100110001";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001100011000";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010110000010";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010010010001";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110011100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010011001101";
        wait for Clk_period; 
        Features_din <= "0000010100011001";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010001100110";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000010011100001";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000010010101101";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000010001110111";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000010010000110";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000010110101011";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010010101010";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000010011110011";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000000100011100";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000010011101001";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001011011100";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010011000011";
        wait for Clk_period; 
        Features_din <= "0000010001100111";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010010001001";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010010101000";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001100010100";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000010110001111";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000010010111010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010010101001";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010110010100";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110011111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010011101110";
        wait for Clk_period; 
        Features_din <= "0000010100011101";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010011100110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010010101000";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010001101001";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000010001101001";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010011001000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010101111100";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010010001110";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010001101010";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010100000101";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000010010010100";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "1111110010101110";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000010010111010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010001010101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001100011001";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000010100000010";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000010001110010";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000010001100001";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010100001010";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000010011100010";
        wait for Clk_period; 
        Features_din <= "0000010101110011";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010010101111";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000010011011010";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010001011100";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010001111011";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010101100010";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010010100110";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111100001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000010101011011";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010010010110";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000010100011110";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000010010100001";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010011111010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010001100001";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010110100100";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010010100110";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001100011101";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010011100111";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010011001110";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001100010011";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000010010110001";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001100011000";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010010101100";
        wait for Clk_period; 
        Features_din <= "0000010011010001";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000010010011100";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010100001001";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010010100011";
        wait for Clk_period; 
        Features_din <= "0000010111110010";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010011010000";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010011110011";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010010010000";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000010110000001";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000010001111011";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110011110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010011100000";
        wait for Clk_period; 
        Features_din <= "0000010101100001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010010111100";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000010001110000";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000010001110000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000010101000111";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010010000010";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010010001000";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001100011100";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001100010100";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001100011010";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010100001111";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "1111111010010110";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000010010111000";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010001101001";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001100001011";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010010000000";
        wait for Clk_period; 
        Features_din <= "0000010010101101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010001110000";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010010001100";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010011001110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000010010111011";
        wait for Clk_period; 
        Features_din <= "0000010101010001";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000010011001100";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010001111000";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001100100011";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010101110100";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000010001110101";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111001101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010010111000";
        wait for Clk_period; 
        Features_din <= "0000010101010110";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010011101100";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010001111000";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010001100101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000010111000100";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010001100100";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010001110100";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001011110000";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010100011110";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001010010011";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000010001111011";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001100101011";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000010100001010";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010001111101";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000010010110110";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000010011000101";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010011000011";
        wait for Clk_period; 
        Features_din <= "0000010110011001";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010001110100";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010010101111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010101010010";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010010000100";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111001001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010011110011";
        wait for Clk_period; 
        Features_din <= "0000010100010010";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010010010001";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000010010100100";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001100010110";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000010010001000";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010010010101";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010110001101";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010010000001";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000010010011001";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010010100111";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001010000110";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000010010111011";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010010010001";
        wait for Clk_period; 
        Features_din <= "0000010001110010";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000010010100101";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000010100011010";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000010010011001";
        wait for Clk_period; 
        Features_din <= "0000010110001000";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010001100011";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010100101100";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010001111101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001100101010";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010101101010";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000010001110000";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110111100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010010100111";
        wait for Clk_period; 
        Features_din <= "0000010100111000";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000010011110011";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000010010110001";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001100011000";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001011110001";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010010000010";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010001111011";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000010110101110";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000010010010011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010010110010";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000010001011011";
        wait for Clk_period; 
        Features_din <= "0000001100011110";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001100011001";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "1111100010010100";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010011100000";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001100010011";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001011111010";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010010010010";
        wait for Clk_period; 
        Features_din <= "0000010011000000";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010010011100";
        wait for Clk_period; 
        Features_din <= "0000010001011100";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000010010100101";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010100000100";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010010100000";
        wait for Clk_period; 
        Features_din <= "0000010110100011";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000010010101110";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010010111110";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010010100100";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001011110011";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010100100100";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010010001011";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110110010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000010100111110";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010010000011";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010001010000";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000010001011100";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000010011000001";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000010001111011";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000010001101111";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010100101010";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001100101011";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000010100000111";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010001111100";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000010001110111";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010011111111";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000010111000100";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001100001110";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000010001111110";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010011111010";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000010010011111";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001011111111";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010001100100";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000010100011101";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110011001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010011000100";
        wait for Clk_period; 
        Features_din <= "0000010100011001";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000010010101100";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010010101101";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001100101011";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010010101001";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000010010010010";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000010110010000";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010010100110";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001100011100";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010011110111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010001111001";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000010011000111";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000010010001100";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000010010011100";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010001100010";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000010010110010";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010100101101";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010001100111";
        wait for Clk_period; 
        Features_din <= "0000010100110101";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001100100011";
        wait for Clk_period; 
        Features_din <= "0000010010011100";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010011110001";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010001100110";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010010110110";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010101011110";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010001110111";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110110010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010010011011";
        wait for Clk_period; 
        Features_din <= "0000010101111000";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010001001101";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010001100011";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010011000110";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010010011110";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000010001110101";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010011010001";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010010010010";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010110010010";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010001100110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010001011010";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001100100100";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010100011111";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001100001101";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010001101111";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001001001101";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000010011011110";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001100110001";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000010010001000";
        wait for Clk_period; 
        Features_din <= "0000010010100000";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010001001101";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010010101110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000011000010000";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010010111010";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000010001001101";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001100100100";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010011010111";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001100100111";
        wait for Clk_period; 
        Features_din <= "0000001100101101";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010101011001";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000010010100000";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001100101000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110000001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010011010010";
        wait for Clk_period; 
        Features_din <= "0000010011100000";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000010011110001";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010001101001";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000010101100010";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000010001100111";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010001111101";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010001011011";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010001100111";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010101000000";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000000001111110";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010010111010";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000010001010000";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000010010101100";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010011000000";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010010101100";
        wait for Clk_period; 
        Features_din <= "0000010101101000";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010010100100";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001100110000";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010001100110";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010010100000";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010110100100";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010001100001";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110100000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010010010110";
        wait for Clk_period; 
        Features_din <= "0000010011110010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010001010000";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000010011110001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010010000010";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000010110101110";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001100011011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010011101011";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "1111100100001010";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010010110001";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010011001101";
        wait for Clk_period; 
        Features_din <= "0000010001110000";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010001100110";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010100001101";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000010001110000";
        wait for Clk_period; 
        Features_din <= "0000010110010011";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000010010101010";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010010101100";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001100010111";
        wait for Clk_period; 
        Features_din <= "0000001100001111";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000010101101011";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010001101010";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001100011000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110011000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010100001000";
        wait for Clk_period; 
        Features_din <= "0000010011000001";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010010110010";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010001100010";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000010100000101";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000010010111000";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010010101100";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010010010011";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000010101010101";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001100100100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001100100011";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010001100001";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000010011110111";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "1111111011110101";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000010011000111";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010001111001";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000010001111101";
        wait for Clk_period; 
        Features_din <= "0000010010001001";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010011000111";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010010010011";
        wait for Clk_period; 
        Features_din <= "0000010111100011";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010011000100";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010010001100";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010001100010";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010101110011";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110011111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000010011111000";
        wait for Clk_period; 
        Features_din <= "0000010100100010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010001111110";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010011010101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000010010000011";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001100100011";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001011110010";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010010010000";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010010000111";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000010111000110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001100001111";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010010111010";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001011101100";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000010011110111";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000010010100101";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000010011100111";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010100100001";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010010000110";
        wait for Clk_period; 
        Features_din <= "0000010110110000";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000010010010000";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010001111001";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010001101110";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010101110000";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000010010000101";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110111111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010011111011";
        wait for Clk_period; 
        Features_din <= "0000010100100011";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000010100011110";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010010011110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010001101010";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000010010100010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000010110011100";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010001111011";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010001101001";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001100101000";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001011111010";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010011110010";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001010011001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000010010111110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001100010000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000010011110011";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010001100101";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000010010000101";
        wait for Clk_period; 
        Features_din <= "0000010110000001";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010010101111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010011101101";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001100000110";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001100010000";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010101001010";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010001100010";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110100111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010001001101";
        wait for Clk_period; 
        Features_din <= "0000010101001101";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000010010100110";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001100001000";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001100100010";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001100001011";
        wait for Clk_period; 
        Features_din <= "0000010100010111";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001011100111";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010001010000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010001010000";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "1111111010111010";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000010010011111";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010010011100";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010011000010";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010010111010";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000010001100101";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010011000000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010011000000";
        wait for Clk_period; 
        Features_din <= "0000010110010110";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010010011101";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010011001000";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000001100001101";
        wait for Clk_period; 
        Features_din <= "0000001100110010";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010101111100";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001100111000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111100110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000010010100100";
        wait for Clk_period; 
        Features_din <= "0000010101000111";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000010010110010";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001100110001";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010010100111";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001100101000";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000010001011100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010010000001";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010110111001";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010001110111";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001100101001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001100001100";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010011101000";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010001110100";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001000101111";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000010011010101";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000010011010110";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010011101001";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000010001110111";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000001100100011";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000010001101001";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010011101111";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001100111000";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000010011000110";
        wait for Clk_period; 
        Features_din <= "0000010110001110";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000010011101111";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010001100100";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000010010011101";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010010000101";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010101011110";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010010010010";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001101100100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010100101011";
        wait for Clk_period; 
        Features_din <= "0000010101001010";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000010100010010";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010010011101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001100000100";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010010000101";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010001100111";
        wait for Clk_period; 
        Features_din <= "0000010010100000";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010001110111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000010101001101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010010010101";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000010001111100";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010100011001";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001100100100";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000010011111001";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010001100001";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001100101010";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000010010010111";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000010011010111";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000010001111000";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010011001110";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000010110010010";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010011001011";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010001110001";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010010111001";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010101110111";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010010010101";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001101101011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000010001010101";
        wait for Clk_period; 
        Features_din <= "0000010101011011";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000010011110010";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010010101100";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001100100011";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010001111011";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010010010001";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000010110001111";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010010100110";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010010100101";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001100101000";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010010100110";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000000101100000";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000010011010101";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000010001111011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001100010110";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000010010011001";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010010101000";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010100000001";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010001011101";
        wait for Clk_period; 
        Features_din <= "0000010110101101";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000010010100011";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010011000100";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001100001001";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010001110100";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010101000011";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010001101010";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111100001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010011101011";
        wait for Clk_period; 
        Features_din <= "0000010110001101";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010010010110";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010100100101";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010010010011";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001100010000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001100100011";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010100110010";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "1111111010111111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000010011001111";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010010010010";
        wait for Clk_period; 
        Features_din <= "0000010010111011";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001100011100";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010001010101";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010011100010";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000010010101010";
        wait for Clk_period; 
        Features_din <= "0000011000101011";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001100101011";
        wait for Clk_period; 
        Features_din <= "0000010010111100";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010010001011";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001100010100";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010110100001";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110100001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000010011010101";
        wait for Clk_period; 
        Features_din <= "0000010101001010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000010010110011";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001100100010";
        wait for Clk_period; 
        Features_din <= "0000010011100001";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010101110011";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010001111000";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010010100000";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001100001110";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010011111011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000010010111010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010010100111";
        wait for Clk_period; 
        Features_din <= "0000010010001010";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001011101000";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000010001001101";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010010111010";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010010111100";
        wait for Clk_period; 
        Features_din <= "0000010111001000";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000010010100110";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000010010011011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010010000000";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001100010011";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010010010111";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010101101100";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010010011010";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001101111011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010010011011";
        wait for Clk_period; 
        Features_din <= "0000010101100010";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000010001100101";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010011000010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000010001101110";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010001100111";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010110001100";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000010001011100";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001100000011";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001100011111";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010011100000";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001100010011";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000010011111000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010010110001";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000001100111000";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000010010101111";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000010001011010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000010001111000";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000010010000001";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010001010000";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010010111010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010011001011";
        wait for Clk_period; 
        Features_din <= "0000010101101011";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010010001101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010010010111";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001100001010";
        wait for Clk_period; 
        Features_din <= "0000001100101011";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010001100011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010101001100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001100100100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111100110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010010101010";
        wait for Clk_period; 
        Features_din <= "0000010110001101";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010001011011";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000010011101111";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000010010000111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010010001011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000010101100111";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010010001000";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010001010000";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000010010000001";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001100110001";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010011111011";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010011111101";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000010010110110";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000010001001101";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000010010000011";
        wait for Clk_period; 
        Features_din <= "0000010010111110";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010001101111";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000010011011101";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010011000011";
        wait for Clk_period; 
        Features_din <= "0000010110010010";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010011100001";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010010101010";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001100011001";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010110011001";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001100011110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110110001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010011010011";
        wait for Clk_period; 
        Features_din <= "0000010100101010";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000010100001001";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001100110000";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010010111110";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000010010110011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010001100011";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001100000101";
        wait for Clk_period; 
        Features_din <= "0000010110001110";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010010011010";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010001100111";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010011011000";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001001101010";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000010100001010";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000010001110001";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000010010100011";
        wait for Clk_period; 
        Features_din <= "0000010010100101";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000010010011001";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000010001100011";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000010010011011";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010011001111";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010010001010";
        wait for Clk_period; 
        Features_din <= "0000010110011100";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010001101110";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000010010100000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001011011000";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001100100110";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010100101111";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010001111110";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110101010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000010100111011";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010001100111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010010100110";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010001100101";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000010110010101";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010001111011";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000010010001101";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001011100110";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001100101000";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010011010100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010010001111";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "1111111011100101";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000010011010110";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000010001001101";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000010011101111";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010001100110";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000010011001001";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010010101100";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000010110001111";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010010001011";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010010100001";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010010011000";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010101010010";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110100101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010010101011";
        wait for Clk_period; 
        Features_din <= "0000010011011111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010011100001";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000010010110000";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000010010101010";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010010010100";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000010110000111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000010001110001";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000010001101001";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010001110100";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001100101011";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001100001001";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001100101000";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010010110001";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000010011100110";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010001001101";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001100100110";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010010000100";
        wait for Clk_period; 
        Features_din <= "0000010001100011";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010010001010";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010011010100";
        wait for Clk_period; 
        Features_din <= "0000010110110100";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001100011000";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001100100010";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000010010010000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010100111100";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010010101011";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111011110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001100010010";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010010110010";
        wait for Clk_period; 
        Features_din <= "0000010100001101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010011010110";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010010100000";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001100011100";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010010011100";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000010101010101";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000010010010001";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010001100111";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010100011001";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "1111111001011010";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000010011001010";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001100001010";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000010001111100";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010010110110";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010011000000";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001100110010";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010010011110";
        wait for Clk_period; 
        Features_din <= "0000010110100000";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001100100110";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010010000011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010010000100";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010010000111";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001100110000";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010111111000";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010010011110";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111110010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010011011100";
        wait for Clk_period; 
        Features_din <= "0000010100111001";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001100101000";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000010011111100";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000010010000001";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010001101111";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010001011100";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000010110111001";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010011010100";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010001101111";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001100110000";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001100010111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010010010011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001010010000";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000010011010100";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000010001101010";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010011000010";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000010010110000";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001100100010";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000010110010101";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010010111000";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010010100100";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010010001111";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010010110011";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110110101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010010000011";
        wait for Clk_period; 
        Features_din <= "0000010011100100";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001100110001";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000010001110111";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010011100100";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000010001011100";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010001001101";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000010110110001";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010010001000";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010001111101";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001011100111";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010011111100";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "1111111111000110";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010011010011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000010010110110";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001100011000";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000010010000100";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010010000011";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010001111110";
        wait for Clk_period; 
        Features_din <= "0000010111000111";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000010001100111";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010011000101";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010001011010";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010001100011";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010100101011";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110101101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010010111010";
        wait for Clk_period; 
        Features_din <= "0000010011011100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010010100101";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000010010100110";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000010001111011";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010011110010";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000010101110000";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000010010101110";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010010000001";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000010011111000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000000010101110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000010010000010";
        wait for Clk_period; 
        Features_din <= "0000010010001011";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010001111000";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010100011011";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000010010101000";
        wait for Clk_period; 
        Features_din <= "0000010110011110";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001100100111";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010010010110";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010010101000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001100011000";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010101101011";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "0000010010000011";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001101111111";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001100110001";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010010011110";
        wait for Clk_period; 
        Features_din <= "0000010100000000";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000010010001111";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010010001101";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010010010010";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010010111111";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001100100110";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010011011110";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010010101110";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001100011110";
        wait for Clk_period; 
        Features_din <= "0000010101110001";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010010001000";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001011111111";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001100110000";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010010000000";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000010011010100";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010001010111";
        wait for Clk_period; 
        Features_din <= "0000001100011101";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010001110100";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000010010100100";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010100000100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001011100111";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010001111101";
        wait for Clk_period; 
        Features_din <= "0000010110100100";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000010010000101";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010001111110";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001100100011";
        wait for Clk_period; 
        Features_din <= "0000001011100101";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010010010010";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010110011001";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010010010100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111010011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010011001101";
        wait for Clk_period; 
        Features_din <= "0000010100000101";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000010001110110";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010001010000";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000010011111101";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010010100010";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001100101101";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010011110110";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000010100011000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001100100100";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010001110111";
        wait for Clk_period; 
        Features_din <= "0000010010000001";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010010011010";
        wait for Clk_period; 
        Features_din <= "0000010001010101";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010011110110";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010010110010";
        wait for Clk_period; 
        Features_din <= "0000010101101101";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000010011000000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010010010011";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010010110010";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001100110001";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001100011010";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010010011110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010110011000";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010011010001";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110011110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010101010010";
        wait for Clk_period; 
        Features_din <= "0000010101000001";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000010100001000";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000010011000010";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010010000110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010001101111";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010100100010";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010001101001";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000010010100001";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010010001100";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001100011000";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001100110010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010010000101";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010011011001";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000010010101011";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000010001011010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000010001010101";
        wait for Clk_period; 
        Features_din <= "0000010011011000";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010001111000";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000010010110001";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001011110010";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010011111000";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001100101011";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010011001011";
        wait for Clk_period; 
        Features_din <= "0000010111011111";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010010101101";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010011000101";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000010010011111";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000010110111001";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010010010011";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001100100110";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001101111011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001100001100";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010010011101";
        wait for Clk_period; 
        Features_din <= "0000010101110101";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010001111101";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000010010011110";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000010010110000";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010001100110";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010001111000";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000010101101000";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010001101111";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010011001111";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010001010101";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001011101111";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010001001101";
        wait for Clk_period; 
        Features_din <= "0000010011011110";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000010001100101";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010010100100";
        wait for Clk_period; 
        Features_din <= "0000010100000111";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000010010100100";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010100001000";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010010100010";
        wait for Clk_period; 
        Features_din <= "0000010110101000";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010010011100";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010011011100";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010101100110";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000010010011001";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110100001";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000010010111101";
        wait for Clk_period; 
        Features_din <= "0000010100000001";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000010001110000";
        wait for Clk_period; 
        Features_din <= "0000010001011011";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010011101101";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010010001010";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010010101001";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010001101110";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000010101011111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001100000111";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010010100001";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000010100000001";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001100110001";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000010010110101";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010010001011";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010011001011";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010010001111";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010010100000";
        wait for Clk_period; 
        Features_din <= "0000010110100001";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000010010101111";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010001111011";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001011111101";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010010101001";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010110110000";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001101101000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010011110011";
        wait for Clk_period; 
        Features_din <= "0000010010110011";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000010001110111";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000010010011000";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010110110011";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010010001101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010001100001";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010001010000";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010101001000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000000001001111";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000010010111101";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001100101000";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010010010100";
        wait for Clk_period; 
        Features_din <= "0000010011100100";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010011010001";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000010001100110";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010101000100";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010010100100";
        wait for Clk_period; 
        Features_din <= "0000010110010011";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000010001110001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010010110011";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000010100001101";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001100100011";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010011010011";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111010010";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010010110001";
        wait for Clk_period; 
        Features_din <= "0000010101111000";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010001111110";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010100010011";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010001111001";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000010110101100";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000010001101010";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010100000000";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "1111111100000111";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001100010110";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000010001110001";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010001101111";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010001100100";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010011100010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000010010010010";
        wait for Clk_period; 
        Features_din <= "0000010111010000";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010011001000";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010011001111";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001100111000";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010100010110";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001100110001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110111101";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010001100010";
        wait for Clk_period; 
        Features_din <= "0000010101100011";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000010001011011";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000010001100101";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000010011010011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000010010001100";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010001100011";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010010101010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010010010101";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010110111110";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010010001011";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010010100110";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010010000110";
        wait for Clk_period; 
        Features_din <= "0000010001010011";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010001011100";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010011011100";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000000110101000";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000010011110100";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001100100011";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010010010010";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010010001101";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000010010100010";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010010100111";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010001110111";
        wait for Clk_period; 
        Features_din <= "0000010111010011";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000010010000100";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010011111001";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010001111011";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001100011110";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010110010111";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010010010100";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001101101100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010011010001";
        wait for Clk_period; 
        Features_din <= "0000010010110101";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000010100000011";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000010001111100";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010010100100";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010001011011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010110000101";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010001111110";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010001100011";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001100011001";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010011100110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001011110001";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000010010111011";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010001111011";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001100110001";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000010010001011";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010010000001";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010001101010";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000010001010000";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001011101100";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010100000000";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010010101011";
        wait for Clk_period; 
        Features_din <= "0000010111000001";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "0000010011011101";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010011001000";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010011001111";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010101110010";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010010000010";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(4, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110100011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010011100001";
        wait for Clk_period; 
        Features_din <= "0000010100000011";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010010000011";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000010011110100";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000010001011100";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000010001110001";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001100110111";
        wait for Clk_period; 
        Features_din <= "0000010101001111";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010001011100";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010001100110";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000010010110000";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000010001011100";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001100111010";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010011110000";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000000011101000";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000010010100100";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000010001100101";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010010110000";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010010000010";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010010100011";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000010100000101";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010010111001";
        wait for Clk_period; 
        Features_din <= "0000010110011100";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000010001101000";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000010011011001";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010011010011";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010101010111";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010010110010";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(3, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110110000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010001111100";
        wait for Clk_period; 
        Features_din <= "0000010101010100";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010001011011";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000010100000101";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000010001111000";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010010000011";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000010110100001";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010000110010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010010010100";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010010011000";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000010011000001";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000000010011111";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000010011001100";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001100101011";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010010100011";
        wait for Clk_period; 
        Features_din <= "0000010001111100";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010010101100";
        wait for Clk_period; 
        Features_din <= "0000010000111111";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000010001100110";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000010001010110";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010001101001";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000010011010100";
        wait for Clk_period; 
        Features_din <= "0000010110000101";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000010010010010";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000010011000111";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001100101000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010101000110";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(2, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110111011";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010001110010";
        wait for Clk_period; 
        Features_din <= "0000010100100111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000010011011000";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010010111111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001100110001";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010010001111";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010110001011";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010001110100";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000010001010000";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010001111101";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010010000010";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010001001000";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000010011111011";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000010000111010";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000010010010011";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010010001000";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010001001110";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010011101100";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010010101010";
        wait for Clk_period; 
        Features_din <= "0000010110011001";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010001100111";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010001110100";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010001100111";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010010100011";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010101101111";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000010010011011";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110010100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010011111110";
        wait for Clk_period; 
        Features_din <= "0000010110000101";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000010001110001";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001011101011";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000010010001000";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001100111000";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010001011101";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010111001111";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000010001100011";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010010011000";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001100010000";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001100000010";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000010001101111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000110011";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "1111110100111110";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000010011101010";
        wait for Clk_period; 
        Features_din <= "0000001100100111";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000010000111011";
        wait for Clk_period; 
        Features_din <= "0000010011110100";
        wait for Clk_period; 
        Features_din <= "0000001100011110";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010010101000";
        wait for Clk_period; 
        Features_din <= "0000010001011100";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000010010101000";
        wait for Clk_period; 
        Features_din <= "0000010000000001";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010100010010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010010101100";
        wait for Clk_period; 
        Features_din <= "0000010100011110";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010001010010";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000010011000010";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000010010111010";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001101001110";
        wait for Clk_period; 
        Features_din <= "0000001100111000";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001100001011";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001100011100";
        wait for Clk_period; 
        Features_din <= "0000001100100001";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010101101000";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010010111110";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(0, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110011000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010011000101";
        wait for Clk_period; 
        Features_din <= "0000010001101111";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010001110000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000010001100101";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001100101000";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001100010111";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000010001101011";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000010101001010";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010000110001";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000010001110100";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001011110101";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001100110000";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000010010010110";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010001011011";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "1111111010100001";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000010010111110";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001101000100";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001100100101";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001100011101";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000010010001110";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010010010001";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000010010110100";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010011111001";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001100110100";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010010110101";
        wait for Clk_period; 
        Features_din <= "0000011000001001";
        wait for Clk_period; 
        Features_din <= "0000001101001010";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001101000110";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010011001110";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010011101010";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001100011000";
        wait for Clk_period; 
        Features_din <= "0000001100110011";
        wait for Clk_period; 
        Features_din <= "0000001100111101";
        wait for Clk_period; 
        Features_din <= "0000001111100011";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001101111010";
        wait for Clk_period; 
        Features_din <= "0000010010000001";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001101001001";
        wait for Clk_period; 
        Features_din <= "0000010101011010";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001100011101";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110001110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001100100000";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000010011000100";
        wait for Clk_period; 
        Features_din <= "0000010011001001";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010010100100";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000010001000111";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000010011110111";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010010000011";
        wait for Clk_period; 
        Features_din <= "0000001100001111";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001100111000";
        wait for Clk_period; 
        Features_din <= "0000001100110000";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000010001011001";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010010111110";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010010000100";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000101010";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010000111000";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000010111011011";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010001011101";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010001110100";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001100101100";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111110110";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000010100010000";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001011011010";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000010011111100";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000010001111100";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000010010001101";
        wait for Clk_period; 
        Features_din <= "0000010011011110";
        wait for Clk_period; 
        Features_din <= "0000001100001001";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010011100101";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000010001100011";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010011001010";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001100111100";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000010010010110";
        wait for Clk_period; 
        Features_din <= "0000011000000000";
        wait for Clk_period; 
        Features_din <= "0000001101101100";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001100010101";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110001001";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010100001111";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000010011101010";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001100111001";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001101000101";
        wait for Clk_period; 
        Features_din <= "0000001100110000";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010110000011";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010001110100";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001101000111";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110111100";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010011000101";
        wait for Clk_period; 
        Features_din <= "0000010100101110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001101101001";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000010000010000";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000010011100111";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101011101";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010001111000";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010000001110";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000010001010100";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010001110101";
        wait for Clk_period; 
        Features_din <= "0000001111010011";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000010001011100";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010001010000";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001101000000";
        wait for Clk_period; 
        Features_din <= "0000010110000000";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000010001011101";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110001101";
        wait for Clk_period; 
        Features_din <= "0000010000010010";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010000101101";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000010001000000";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111001010";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010010100101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000010000100011";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000000110011001";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000010011100001";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001100111111";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000010010001000";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010000100111";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000010011000101";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001101110110";
        wait for Clk_period; 
        Features_din <= "0000010010100001";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001100100111";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000010010101000";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000010001110001";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001101010101";
        wait for Clk_period; 
        Features_din <= "0000010000111101";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010010111011";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001100101110";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000010010110111";
        wait for Clk_period; 
        Features_din <= "0000010110100101";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010011000110";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010100110100";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001100111000";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010001101111";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111011111";
        wait for Clk_period; 
        Features_din <= "0000001100110000";
        wait for Clk_period; 
        Features_din <= "0000001101100100";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000010001100110";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010101111001";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000010000100101";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001111010110";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000010010101111";
        wait for Clk_period; 
        Features_din <= "0000010100110000";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000010000010101";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001101001000";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000010001011111";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000010010110001";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000010000011000";
        wait for Clk_period; 
        Features_din <= "0000001100100110";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000010001110010";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000010000011011";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000010010111101";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000010001011000";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000010110101101";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000010001001111";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010011001011";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110001011";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010000111100";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001101010000";
        wait for Clk_period; 
        Features_din <= "0000001111101111";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001100100011";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000010000000110";
        wait for Clk_period; 
        Features_din <= "0000001111111100";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010011100111";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000010000101001";
        wait for Clk_period; 
        Features_din <= "0000000010001111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000010011111111";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010000110111";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001101010011";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010000100110";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001100001000";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111111010";
        wait for Clk_period; 
        Features_din <= "0000001101011100";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000010001111010";
        wait for Clk_period; 
        Features_din <= "0000001101100110";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000010011011100";
        wait for Clk_period; 
        Features_din <= "0000010000001111";
        wait for Clk_period; 
        Features_din <= "0000010001100000";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001101100001";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010010100101";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010010010011";
        wait for Clk_period; 
        Features_din <= "0000010110011111";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001101000011";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000010010001100";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000010010100111";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001101111011";
        wait for Clk_period; 
        Features_din <= "0000010001111111";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000010000001001";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001101010111";
        wait for Clk_period; 
        Features_din <= "0000001111000110";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010110110111";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000010010000110";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001100011001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110101000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001111000000";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111111011";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010011101110";
        wait for Clk_period; 
        Features_din <= "0000010010111010";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001101100101";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001111010101";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010000000101";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000010001011010";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000010011101000";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010010100001";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111111000";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001111011110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001100111011";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010000010001";
        wait for Clk_period; 
        Features_din <= "0000010000100010";
        wait for Clk_period; 
        Features_din <= "0000001110110010";
        wait for Clk_period; 
        Features_din <= "0000001110011001";
        wait for Clk_period; 
        Features_din <= "0000010001111110";
        wait for Clk_period; 
        Features_din <= "0000001110110110";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001110011111";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000010000101111";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001110010010";
        wait for Clk_period; 
        Features_din <= "0000010110000011";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010001000100";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010000111110";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000010010010100";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000010001111001";
        wait for Clk_period; 
        Features_din <= "0000001111111111";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001101110000";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000010000001010";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001110011101";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000010000011010";
        wait for Clk_period; 
        Features_din <= "0000001100111110";
        wait for Clk_period; 
        Features_din <= "0000001111010100";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        Features_din <= "0000001101101111";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001111100010";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010000000111";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111100101";
        wait for Clk_period; 
        Features_din <= "0000001111011000";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000010010011011";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000010000100001";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000010001010001";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001100010000";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111000111";
        wait for Clk_period; 
        Features_din <= "0000010000101100";
        wait for Clk_period; 
        Features_din <= "0000010011010010";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110001010";
        wait for Clk_period; 
        Features_din <= "0000001111100000";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001101100111";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000010000011110";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001100110101";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010000110000";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010000011100";
        wait for Clk_period; 
        Features_din <= "0000001111110101";
        wait for Clk_period; 
        Features_din <= "0000001101110010";
        wait for Clk_period; 
        Features_din <= "0000010010001101";
        wait for Clk_period; 
        Features_din <= "0000010011000100";
        wait for Clk_period; 
        Features_din <= "0000001110100100";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000010001110111";
        wait for Clk_period; 
        Features_din <= "0000010000000010";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000010000101011";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010010100101";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000010000011101";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110010101";
        wait for Clk_period; 
        Features_din <= "0000001101011111";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001101011010";
        wait for Clk_period; 
        Features_din <= "0000010000101110";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001101111110";
        wait for Clk_period; 
        Features_din <= "0000010010110101";
        wait for Clk_period; 
        Features_din <= "0000001110010000";
        wait for Clk_period; 
        Features_din <= "0000001110101011";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000001101010001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000010001101001";
        wait for Clk_period; 
        Features_din <= "0000010110000011";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001111110111";
        wait for Clk_period; 
        Features_din <= "0000001100110110";
        wait for Clk_period; 
        Features_din <= "0000001110101111";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000010001000001";
        wait for Clk_period; 
        Features_din <= "0000001110101010";
        wait for Clk_period; 
        Features_din <= "0000001110000111";
        wait for Clk_period; 
        Features_din <= "0000001101111000";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000010001100001";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000010010111010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000001111001100";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001110101000";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001101110100";
        wait for Clk_period; 
        Features_din <= "0000010011010110";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001111101110";
        wait for Clk_period; 
        Features_din <= "0000001101101110";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000001111010111";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000010001101110";
        wait for Clk_period; 
        Features_din <= "0000001110000001";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000010110100111";
        wait for Clk_period; 
        Features_din <= "0000001111101011";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000001111110100";
        wait for Clk_period; 
        Features_din <= "0000001101010010";
        wait for Clk_period; 
        Features_din <= "0000001101011001";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
        class_label <= std_logic_vector(to_unsigned(1, class_label'length));
        
        -- Load and valid features flags
        Load_features <= '1';
        Valid_feature <= '1';
        
        Features_din <= "0000001110101000";
        wait for Clk_period;

        -- Reset load flag
        Load_features <= '0';
        
        Features_din <= "0000001111101000";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000010000100000";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110000010";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010010101010";
        wait for Clk_period; 
        Features_din <= "0000010101110001";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000010000100100";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111100001";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110001000";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000010001001011";
        wait for Clk_period; 
        Features_din <= "0000001110001100";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001101100000";
        wait for Clk_period; 
        Features_din <= "0000010001001100";
        wait for Clk_period; 
        Features_din <= "0000001111000100";
        wait for Clk_period; 
        Features_din <= "0000010001000110";
        wait for Clk_period; 
        Features_din <= "0000010001100100";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000010001011110";
        wait for Clk_period; 
        Features_din <= "0000001110101100";
        wait for Clk_period; 
        Features_din <= "0000001110011110";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010011110100";
        wait for Clk_period; 
        Features_din <= "0000001111000001";
        wait for Clk_period; 
        Features_din <= "0000010000011111";
        wait for Clk_period; 
        Features_din <= "0000001101001111";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111110011";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000010000001100";
        wait for Clk_period; 
        Features_din <= "0000001011111000";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000010000110110";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000001101010100";
        wait for Clk_period; 
        Features_din <= "0000010001110011";
        wait for Clk_period; 
        Features_din <= "0000001111000011";
        wait for Clk_period; 
        Features_din <= "0000001101001011";
        wait for Clk_period; 
        Features_din <= "0000001101000001";
        wait for Clk_period; 
        Features_din <= "0000010010101011";
        wait for Clk_period; 
        Features_din <= "0000001111011001";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000010000010100";
        wait for Clk_period; 
        Features_din <= "0000001101111111";
        wait for Clk_period; 
        Features_din <= "0000010110010100";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001110110011";
        wait for Clk_period; 
        Features_din <= "0000001111100111";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001111110010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000010001110010";
        wait for Clk_period; 
        Features_din <= "0000001110111000";
        wait for Clk_period; 
        Features_din <= "0000010010001011";
        wait for Clk_period; 
        Features_din <= "0000001111011011";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111100110";
        wait for Clk_period; 
        Features_din <= "0000001101110111";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001101101101";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110010111";
        wait for Clk_period; 
        Features_din <= "0000001101011110";
        wait for Clk_period; 
        Features_din <= "0000001111110001";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000010001000011";
        wait for Clk_period; 
        Features_din <= "0000010000101000";
        wait for Clk_period; 
        Features_din <= "0000001110111100";
        wait for Clk_period; 
        Features_din <= "0000001110000101";
        wait for Clk_period; 
        Features_din <= "0000001111101101";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001110011010";
        wait for Clk_period; 
        Features_din <= "0000010000000000";
        wait for Clk_period; 
        Features_din <= "0000001100100100";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101111100";
        wait for Clk_period; 
        Features_din <= "0000001101000010";
        wait for Clk_period; 
        Features_din <= "0000001101100011";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111011101";
        wait for Clk_period; 
        Features_din <= "0000001100100110";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110000110";
        wait for Clk_period; 
        Features_din <= "0000010001001001";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000010000011001";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111001111";
        wait for Clk_period; 
        Features_din <= "0000001111100100";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000001110100111";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000010000001011";
        wait for Clk_period; 
        Features_din <= "0000001101110101";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001111101001";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000001111001011";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000010011000001";
        wait for Clk_period; 
        Features_din <= "0000001110110100";
        wait for Clk_period; 
        Features_din <= "0000001101111101";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001111111101";
        wait for Clk_period; 
        Features_din <= "0000001111110000";
        wait for Clk_period; 
        Features_din <= "0000001110110001";
        wait for Clk_period; 
        Features_din <= "0000010010001010";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001110110111";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110101110";
        wait for Clk_period; 
        Features_din <= "0000001111001110";
        wait for Clk_period; 
        Features_din <= "0000001000111011";
        wait for Clk_period; 
        Features_din <= "0000001111011100";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000010001000101";
        wait for Clk_period; 
        Features_din <= "0000010011001110";
        wait for Clk_period; 
        Features_din <= "0000001110110000";
        wait for Clk_period; 
        Features_din <= "0000001110111011";
        wait for Clk_period; 
        Features_din <= "0000010001011011";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000010000111001";
        wait for Clk_period; 
        Features_din <= "0000001101010110";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000010000001000";
        wait for Clk_period; 
        Features_din <= "0000010001101100";
        wait for Clk_period; 
        Features_din <= "0000001111000101";
        wait for Clk_period; 
        Features_din <= "0000001111010001";
        wait for Clk_period; 
        Features_din <= "0000001111101010";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110000100";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001101101000";
        wait for Clk_period; 
        Features_din <= "0000010001100010";
        wait for Clk_period; 
        Features_din <= "0000010010110010";
        wait for Clk_period; 
        Features_din <= "0000001100011000";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111010110";
        wait for Clk_period; 
        Features_din <= "0000010001001010";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000001101011011";
        wait for Clk_period; 
        Features_din <= "0000010000010110";
        wait for Clk_period; 
        Features_din <= "0000001110011100";
        wait for Clk_period; 
        Features_din <= "0000001111010010";
        wait for Clk_period; 
        Features_din <= "0000001110000011";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000010011000110";
        wait for Clk_period; 
        Features_din <= "0000010000010111";
        wait for Clk_period; 
        Features_din <= "0000010001101101";
        wait for Clk_period; 
        Features_din <= "0000001111001101";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110100101";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000001110100000";
        wait for Clk_period; 
        Features_din <= "0000001100011111";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000010000110100";
        wait for Clk_period; 
        Features_din <= "0000010000001101";
        wait for Clk_period; 
        Features_din <= "0000001110010110";
        wait for Clk_period; 
        Features_din <= "0000010010001001";
        wait for Clk_period; 
        Features_din <= "0000001110111101";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110101101";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001110010001";
        wait for Clk_period; 
        Features_din <= "0000010000000100";
        wait for Clk_period; 
        Features_din <= "0000010010010100";
        wait for Clk_period; 
        Features_din <= "0000010110010100";
        wait for Clk_period; 
        Features_din <= "0000001110010100";
        wait for Clk_period; 
        Features_din <= "0000001110100011";
        wait for Clk_period; 
        Features_din <= "0000001110111010";
        wait for Clk_period; 
        Features_din <= "0000001111111110";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110110101";
        wait for Clk_period; 
        Features_din <= "0000001101110001";
        wait for Clk_period; 
        Features_din <= "0000001101101010";
        wait for Clk_period; 
        Features_din <= "0000010000010011";
        wait for Clk_period; 
        Features_din <= "0000001110100110";
        wait for Clk_period; 
        Features_din <= "0000001101101011";
        wait for Clk_period; 
        Features_din <= "0000001101100010";
        wait for Clk_period; 
        Features_din <= "0000001101001100";
        wait for Clk_period; 
        Features_din <= "0000010010010111";
        wait for Clk_period; 
        Features_din <= "0000001101111001";
        wait for Clk_period; 
        Features_din <= "0000010010111000";
        wait for Clk_period; 
        Features_din <= "0000001110101001";
        wait for Clk_period; 
        Features_din <= "0000001100011011";
        wait for Clk_period; 
        Features_din <= "0000001111101100";
        wait for Clk_period; 
        Features_din <= "0000001110001111";
        wait for Clk_period; 
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        Features_din <= "0000001110000000";
        wait for Clk_period; 
        Features_din <= "0000001110011011";
        wait for Clk_period; 
        Features_din <= "0000010011000111";
        wait for Clk_period; 
        Features_din <= "0000001110001110";
        wait for Clk_period; 
        Features_din <= "0000001111111001";
        wait for Clk_period; 
        Features_din <= "0000001110100001";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110111110";
        wait for Clk_period; 
        Features_din <= "0000001111000010";
        wait for Clk_period; 
        Features_din <= "0000001100101111";
        wait for Clk_period; 
        Features_din <= "0000001100001101";
        wait for Clk_period; 
        Features_din <= "0000001101110011";
        wait for Clk_period; 
        Features_din <= "0000001111001001";
        wait for Clk_period; 
        Features_din <= "0000010000110101";
        wait for Clk_period; 
        Features_din <= "0000001110010011";
        wait for Clk_period; 
        Features_din <= "0000001110100010";
        wait for Clk_period; 
        Features_din <= "0000010001000010";
        wait for Clk_period; 
        Features_din <= "0000001110111111";
        wait for Clk_period; 
        Features_din <= "0000001110011000";
        wait for Clk_period; 
        Features_din <= "0000010100110100";
        wait for Clk_period; 
        Features_din <= "0000010000000011";
        wait for Clk_period; 
        Features_din <= "0000001111010000";
        wait for Clk_period; 
        Features_din <= "0000001110111001";
        wait for Clk_period; 
        Features_din <= "0000010001111000";
        wait for Clk_period; 
        Features_din <= "0000001111011010";
        wait for Clk_period; 
        Features_din <= "0000001101001101";
        wait for Clk_period; 
        Features_din <= "0000001101011000";
        wait for Clk_period; 
        

        last_feature <= '1';
        pc_count     <= '1'; -- count pixel
        Features_din <= "0000001111001000";
        wait for Clk_period; 
        
        

        -- Reset count, last and valid flags
        pc_count      <= '0';
        Last_feature  <= '0';
        Valid_feature <= '0';
        
        -- Wait until inference is complete
        wait until Finish = '1';
        
        wait for Clk_period * 1/2;
        
        if Dout = class_label then
            hc_count <= '1';
        end if;
        
        wait for Clk_period;
        hc_count <= '0';
        
        
            wait;
    end process;
end;
